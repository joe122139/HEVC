`timescale 1ns/1ps
module intra_pseudoAddr(
	mode,			//i
	X,				//i
	Y,
	pseuAdr
	,preStage		//input    0:pre0;  1:pre1;    4: calculation stage
	,tuSize			//input
);

	
	parameter AW = 3;
	
	input [5:0] mode;
	input [2:0] X;
	input [2:0] Y;
	input [3:0] preStage;   // 0:pre0;  1:pre1;    4: calculation stage
	input [2:0] tuSize;
	
	output reg [AW*8-1:0]   pseuAdr;
	 
	reg [AW-1:0] adrVal [7:0];			// AW * 4;	


	
/*for debug*/
  reg [5:0] r_mode;
	always @(*) begin
		r_mode <= mode;
	end
/*for debug*/

	generate
	  genvar i;
	  for(i=0;i<8;i=i+1) begin:xi
	    always @(*) begin
		    pseuAdr [AW*8-1-AW*i: AW*7-AW*i] = adrVal[i];
	    end
	  end
	endgenerate


always @(*) begin
case(preStage)
4'd0: begin 
	if( mode!=6'd1 && tuSize== 3'd5)		//planar + angular
		begin  adrVal[0]= 3 ; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]=  2 ;  end		//ab [7]  le [0] 	ab,le:63
	else if( mode==0 && tuSize== 3'd4)		//planar, PU16
		begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;  end		//ab[2-4] ab 11-17              (//le [5-3]	  le 11-17)
  else if (mode==6'd1) 
		begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;  end			//ab  0-15
	else 
		begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;  end
 end
4'd1: begin 
	if( mode!=6'd1 && tuSize== 6'd5)		//planar + angular
		begin  adrVal[0]=  1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]=  0;  end		//left　31, ab 31	
	else if (mode==6'd1) 
		begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]=  0; adrVal[5]=  0; adrVal[6]= 0 ; adrVal[7]= 0 ;  end		//ab  16-31
	else 
		begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;  end
	end
	
4'd2: begin 
	if( mode!=6'd1 && tuSize== 6'd5)		//planar + angular
		begin  adrVal[0]=  1; adrVal[1]=  1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]=  3;  end		//left [1] [0] [7]		le:27-33
	else if (mode==6'd1) 
		begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]=  1; adrVal[5]=  1; adrVal[6]= 1 ; adrVal[7]=  1 ;  end		//le  0-15
	else 
		begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;  end
	end
	
4'd3: begin
	if( mode!=6'd1 && tuSize== 6'd5)		//planar + angular
		begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;  end		//above [6] [7] [0]		ab:27-33
	else if (mode==6'd1) 
		begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]=  7; adrVal[5]=  7; adrVal[6]= 7 ; adrVal[7]=  7 ;  end		//le  16-31
	else 
		begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;  end
 end
4'd4: begin
	if (mode==6'd1) 
		begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]=  7; adrVal[5]=  7; adrVal[6]= 7 ; adrVal[7]=  7 ;  end		//ab  32-47
	else 
		begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;  end
 end 
4'd5: begin
	if (mode==6'd1) 
		begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]=  2; adrVal[5]=  2; adrVal[6]= 2 ; adrVal[7]=  2 ;  end		//ab  48-63
	else 
		begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;  end
 end 
4'd6: begin
	if (mode==6'd1) 
		begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]=  3; adrVal[5]=  3; adrVal[6]= 3 ; adrVal[7]=  3 ;  end		//le  32-47
	else 
		begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;  end
 end 
4'd7: begin
	if (mode==6'd1) 
		begin  adrVal[0]= 3; adrVal[1]= 3; adrVal[2]= 3; adrVal[3]= 3; adrVal[4]=  7; adrVal[5]=  7; adrVal[6]= 7 ; adrVal[7]=  7 ;  end		//le  48-63
	else 
		begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;  end
 end  
default: begin
 case({mode,1'b0,X,1'b0,Y})
14'h 000: 
			if(tuSize== 3'd2)	begin		
				adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;		end
			else				begin
			  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;    //0,1,2,3,-1,-1,-1,-1,
		end
14'h 001: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,-1,-1,-1,-1,
14'h 002: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,-1,-1,-1,-1,
14'h 003: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,-1,-1,-1,-1,
14'h 004: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,-1,-1,-1,-1,
14'h 005: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,-1,-1,-1,-1,
14'h 006: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,-1,-1,-1,-1,
14'h 007: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,-1,-1,-1,-1,
14'h 010: if(tuSize==3'd3)
		begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //-1,-1,-1,-1,0,1,2,3
		else
			begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,-1,-1,-1,-1,
14'h 011: if(tuSize==3'd3) 
			begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,4,5,6,7,
		else
			begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,-1,-1,-1,-1,
14'h 012: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,-1,-1,-1,-1,
14'h 013: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,-1,-1,-1,-1,
14'h 014: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,-1,-1,-1,-1,
14'h 015: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,-1,-1,-1,-1,
14'h 016: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,-1,-1,-1,-1,
14'h 017: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,-1,-1,-1,-1,
14'h 020: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h 021: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h 022: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h 023: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h 024: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h 025: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h 026: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h 027: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h 030:   
    if(tuSize==3'd4)
      begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //-1,-1,-1,-1,0,1,2,3,
    else 
      begin adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
  
14'h 031: 
	if(tuSize==3'd4)
      begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //-1,-1,-1,-1,4,5,6,7,
    else 
	begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,

14'h 032: 
	if(tuSize==3'd4)
      begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //-1,-1,-1,-1,8,9,10,11,
    else 
	  begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,

14'h 033: 
	if(tuSize==3'd4)
      begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //-1,-1,-1,-1,12,13,14,15,
	else
	  begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h 034: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h 035: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h 036: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h 037: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h 040: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h 041: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h 042: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h 043: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h 044: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h 045: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h 046: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h 047: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h 050: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h 051: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h 052: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h 053: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h 054: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h 055: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h 056: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h 057: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h 060: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,-1,-1,-1,-1,
14'h 061: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,-1,-1,-1,-1,
14'h 062: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,-1,-1,-1,-1,
14'h 063: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,-1,-1,-1,-1,
14'h 064: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,-1,-1,-1,-1,
14'h 065: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,-1,-1,-1,-1,
14'h 066: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,-1,-1,-1,-1,
14'h 067: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,-1,-1,-1,-1,
14'h 070: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //-1,-1,-1,-1,0,1,2,3,
14'h 071: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //-1,-1,-1,-1,4,5,6,7,
14'h 072: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //-1,-1,-1,-1,8,9,10,11,
14'h 073: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //-1,-1,-1,-1,12,13,14,15,
14'h 074: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //-1,-1,-1,-1,16,17,18,19,
14'h 075: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //-1,-1,-1,-1,20,21,22,23,
14'h 076: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //-1,-1,-1,-1,24,25,26,27,
14'h 077: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //-1,-1,-1,-1,28,29,30,31,
14'h 100: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,0,1,2,3,
14'h 101: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,6,7,
14'h 102: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //0,1,2,3,8,9,10,11,
14'h 103: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,12,13,14,15,
14'h 104: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,16,17,18,19,
14'h 105: begin  adrVal[0]= 0; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,20,21,22,23,
14'h 106: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,24,25,26,27,
14'h 107: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //0,1,2,3,28,29,30,31,
14'h 110: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,0,1,2,3,
14'h 111: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,4,5,6,7,
14'h 112: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //4,5,6,7,8,9,10,11,
14'h 113: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,12,13,14,15,
14'h 114: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,16,17,18,19,
14'h 115: begin  adrVal[0]= 0; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,20,21,22,23,
14'h 116: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,24,25,26,27,
14'h 117: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //4,5,6,7,28,29,30,31,
14'h 120: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //8,9,10,11,0,1,2,3,
14'h 121: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //8,9,10,11,4,5,6,7,
14'h 122: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,8,9,10,11,
14'h 123: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,15,
14'h 124: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,16,17,18,19,
14'h 125: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,20,21,22,23,
14'h 126: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,24,25,26,27,
14'h 127: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //8,9,10,11,28,29,30,31,
14'h 130: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //12,13,14,15,0,1,2,3,
14'h 131: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //12,13,14,15,4,5,6,7,
14'h 132: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //12,13,14,15,8,9,10,11,
14'h 133: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //12,13,14,15,12,13,14,15,
14'h 134: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,19,
14'h 135: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,20,21,22,23,
14'h 136: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,24,25,26,27,
14'h 137: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //12,13,14,15,28,29,30,31,
14'h 140: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 1; adrVal[7]= 1;   end //16,17,18,19,0,1,2,3,
14'h 141: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //16,17,18,19,4,5,6,7,
14'h 142: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //16,17,18,19,8,9,10,11,
14'h 143: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,12,13,14,15,
14'h 144: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,16,17,18,19,
14'h 145: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,23,
14'h 146: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,24,25,26,27,
14'h 147: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 3;   end //16,17,18,19,28,29,30,31,
14'h 150: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 1; adrVal[7]= 1;   end //20,21,22,23,0,1,2,3,
14'h 151: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //20,21,22,23,4,5,6,7,
14'h 152: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //20,21,22,23,8,9,10,11,
14'h 153: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,12,13,14,15,
14'h 154: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,16,17,18,19,
14'h 155: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,20,21,22,23,
14'h 156: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,26,27,
14'h 157: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 3;   end //20,21,22,23,28,29,30,31,
14'h 160: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 1; adrVal[7]= 1;   end //24,25,26,27,0,1,2,3,
14'h 161: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //24,25,26,27,4,5,6,7,
14'h 162: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 0;   end //24,25,26,27,8,9,10,11,
14'h 163: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,12,13,14,15,
14'h 164: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,16,17,18,19,
14'h 165: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,20,21,22,23,
14'h 166: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,24,25,26,27,
14'h 167: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 3;   end //24,25,26,27,28,29,30,31,
14'h 170: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //28,29,30,31,0,1,2,3,
14'h 171: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //28,29,30,31,4,5,6,7,
14'h 172: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 0;   end //28,29,30,31,8,9,10,11,
14'h 173: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,12,13,14,15,
14'h 174: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,16,17,18,19,
14'h 175: begin  adrVal[0]= 2; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,20,21,22,23,
14'h 176: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,24,25,26,27,
14'h 177: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 3;   end //28,29,30,31,28,29,30,31,
14'h 200: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,7,8,
14'h 201: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,11,12,
14'h 202: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,16,
14'h 203: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,20,
14'h 204: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,24,
14'h 205: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,28,
14'h 206: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //25,26,27,28,29,30,31,32,
14'h 207: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //29,30,31,32,33,34,35,36,
14'h 210: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,11,12,
14'h 211: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,16,
14'h 212: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,20,
14'h 213: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,24,
14'h 214: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,28,
14'h 215: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //25,26,27,28,29,30,31,32,
14'h 216: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //29,30,31,32,33,34,35,36,
14'h 217: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //33,34,35,36,37,38,39,40,
14'h 220: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,16,
14'h 221: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,20,
14'h 222: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,24,
14'h 223: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,28,
14'h 224: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //25,26,27,28,29,30,31,32,
14'h 225: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //29,30,31,32,33,34,35,36,
14'h 226: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //33,34,35,36,37,38,39,40,
14'h 227: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //37,38,39,40,41,42,43,44,
14'h 230: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,20,
14'h 231: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,24,
14'h 232: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,28,
14'h 233: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //25,26,27,28,29,30,31,32,
14'h 234: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //29,30,31,32,33,34,35,36,
14'h 235: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //33,34,35,36,37,38,39,40,
14'h 236: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //37,38,39,40,41,42,43,44,
14'h 237: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,48,
14'h 240: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,24,
14'h 241: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,28,
14'h 242: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //25,26,27,28,29,30,31,32,
14'h 243: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //29,30,31,32,33,34,35,36,
14'h 244: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //33,34,35,36,37,38,39,40,
14'h 245: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //37,38,39,40,41,42,43,44,
14'h 246: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,48,
14'h 247: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 3; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //45,46,47,48,49,50,51,52,
14'h 250: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,28,
14'h 251: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //25,26,27,28,29,30,31,32,
14'h 252: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //29,30,31,32,33,34,35,36,
14'h 253: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //33,34,35,36,37,38,39,40,
14'h 254: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //37,38,39,40,41,42,43,44,
14'h 255: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,48,
14'h 256: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 3; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //45,46,47,48,49,50,51,52,
14'h 257: begin  adrVal[0]= 7; adrVal[1]= 3; adrVal[2]= 3; adrVal[3]= 3; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //49,50,51,52,53,54,55,56,
14'h 260: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //25,26,27,28,29,30,31,32,
14'h 261: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //29,30,31,32,33,34,35,36,
14'h 262: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //33,34,35,36,37,38,39,40,
14'h 263: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //37,38,39,40,41,42,43,44,
14'h 264: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,48,
14'h 265: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 3; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //45,46,47,48,49,50,51,52,
14'h 266: begin  adrVal[0]= 7; adrVal[1]= 3; adrVal[2]= 3; adrVal[3]= 3; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //49,50,51,52,53,54,55,56,
14'h 267: begin  adrVal[0]= 3; adrVal[1]= 3; adrVal[2]= 3; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //53,54,55,56,57,58,59,60,
14'h 270: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //29,30,31,32,33,34,35,36,
14'h 271: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //33,34,35,36,37,38,39,40,
14'h 272: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //37,38,39,40,41,42,43,44,
14'h 273: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,48,
14'h 274: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 3; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //45,46,47,48,49,50,51,52,
14'h 275: begin  adrVal[0]= 7; adrVal[1]= 3; adrVal[2]= 3; adrVal[3]= 3; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //49,50,51,52,53,54,55,56,
14'h 276: begin  adrVal[0]= 3; adrVal[1]= 3; adrVal[2]= 3; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //53,54,55,56,57,58,59,60,
14'h 277: begin  adrVal[0]= 3; adrVal[1]= 3; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 5;   end //57,58,59,60,61,62,63,64,
14'h 300: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,6,7,
14'h 301: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,10,11,
14'h 302: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,13,14,
14'h 303: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,17,
14'h 304: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,20,
14'h 305: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,24,
14'h 306: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,26,27,
14'h 307: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,29,30,
14'h 310: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,10,11,
14'h 311: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,14,15,
14'h 312: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,18,
14'h 313: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,21,
14'h 314: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,24,
14'h 315: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,28,
14'h 316: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //24,25,26,27,28,29,30,31,
14'h 317: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,32,33,34,
14'h 320: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,14,15,
14'h 321: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,19,
14'h 322: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,22,
14'h 323: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,24,25,
14'h 324: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,28,
14'h 325: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //25,26,27,28,29,30,31,32,
14'h 326: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //28,29,30,31,32,33,34,35,
14'h 327: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //31,32,33,34,35,36,37,38,
14'h 330: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,19,
14'h 331: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,23,
14'h 332: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,25,26,
14'h 333: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,27,28,29,
14'h 334: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //25,26,27,28,29,30,31,32,
14'h 335: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //29,30,31,32,33,34,35,36,
14'h 336: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //32,33,34,35,36,37,38,39,
14'h 337: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //35,36,37,38,39,40,41,42,
14'h 340: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,23,
14'h 341: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,26,27,
14'h 342: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,29,30,
14'h 343: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //26,27,28,29,30,31,32,33,
14'h 344: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //29,30,31,32,33,34,35,36,
14'h 345: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //33,34,35,36,37,38,39,40,
14'h 346: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //36,37,38,39,40,41,42,43,
14'h 347: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //39,40,41,42,43,44,45,46,
14'h 350: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,26,27,
14'h 351: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //24,25,26,27,28,29,30,31,
14'h 352: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,32,33,34,
14'h 353: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //30,31,32,33,34,35,36,37,
14'h 354: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //33,34,35,36,37,38,39,40,
14'h 355: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //37,38,39,40,41,42,43,44,
14'h 356: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //40,41,42,43,44,45,46,47,
14'h 357: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 7; adrVal[7]= 7;   end //43,44,45,46,47,48,49,50,
14'h 360: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //24,25,26,27,28,29,30,31,
14'h 361: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //28,29,30,31,32,33,34,35,
14'h 362: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //31,32,33,34,35,36,37,38,
14'h 363: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //34,35,36,37,38,39,40,41,
14'h 364: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //37,38,39,40,41,42,43,44,
14'h 365: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,48,
14'h 366: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 3; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 7; adrVal[7]= 7;   end //44,45,46,47,48,49,50,51,
14'h 367: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 3; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //47,48,49,50,51,52,53,54,
14'h 370: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //28,29,30,31,32,33,34,35,
14'h 371: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //32,33,34,35,36,37,38,39,
14'h 372: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //35,36,37,38,39,40,41,42,
14'h 373: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //38,39,40,41,42,43,44,45,
14'h 374: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,48,
14'h 375: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 3; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //45,46,47,48,49,50,51,52,
14'h 376: begin  adrVal[0]= 7; adrVal[1]= 3; adrVal[2]= 3; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //48,49,50,51,52,53,54,55,
14'h 377: begin  adrVal[0]= 7; adrVal[1]= 3; adrVal[2]= 3; adrVal[3]= 3; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //51,52,53,54,55,56,57,58,
14'h 400: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,6,-1,
14'h 401: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,9,-1,
14'h 402: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h 403: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h 404: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h 405: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h 406: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h 407: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h 410: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,10,-1,
14'h 411: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h 412: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h 413: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h 414: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h 415: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h 416: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h 417: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,29,-1,
14'h 420: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h 421: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h 422: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h 423: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h 424: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h 425: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,-1,
14'h 426: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,30,-1,
14'h 427: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,32,33,-1,
14'h 430: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h 431: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h 432: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h 433: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h 434: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,29,-1,
14'h 435: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //25,26,27,28,29,30,31,-1,
14'h 436: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,34,-1,
14'h 437: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //31,32,33,34,35,36,37,-1,
14'h 440: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h 441: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h 442: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,-1,
14'h 443: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,30,-1,
14'h 444: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,32,33,-1,
14'h 445: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //29,30,31,32,33,34,35,-1,
14'h 446: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //32,33,34,35,36,37,38,-1,
14'h 447: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //35,36,37,38,39,40,41,-1,
14'h 450: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h 451: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,29,-1,
14'h 452: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //25,26,27,28,29,30,31,-1,
14'h 453: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,34,-1,
14'h 454: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //31,32,33,34,35,36,37,-1,
14'h 455: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //33,34,35,36,37,38,39,-1,
14'h 456: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //36,37,38,39,40,41,42,-1,
14'h 457: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //39,40,41,42,43,44,45,-1,
14'h 460: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,30,-1,
14'h 461: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,32,33,-1,
14'h 462: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //29,30,31,32,33,34,35,-1,
14'h 463: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //32,33,34,35,36,37,38,-1,
14'h 464: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //35,36,37,38,39,40,41,-1,
14'h 465: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //37,38,39,40,41,42,43,-1,
14'h 466: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //40,41,42,43,44,45,46,-1,
14'h 467: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 7; adrVal[7]= 7;   end //43,44,45,46,47,48,49,-1,
14'h 470: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,34,-1,
14'h 471: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //31,32,33,34,35,36,37,-1,
14'h 472: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //33,34,35,36,37,38,39,-1,
14'h 473: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //36,37,38,39,40,41,42,-1,
14'h 474: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //39,40,41,42,43,44,45,-1,
14'h 475: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,-1,
14'h 476: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 7; adrVal[7]= 7;   end //44,45,46,47,48,49,50,-1,
14'h 477: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 3; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //47,48,49,50,51,52,53,-1,
14'h 500: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,6,-1,
14'h 501: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,7,8,-1,
14'h 502: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,10,-1,
14'h 503: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,11,12,-1,
14'h 504: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h 505: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h 506: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h 507: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h 510: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,10,-1,
14'h 511: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,11,12,-1,
14'h 512: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h 513: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h 514: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h 515: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h 516: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h 517: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h 520: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h 521: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h 522: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h 523: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h 524: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h 525: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h 526: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,-1,
14'h 527: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,29,-1,
14'h 530: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h 531: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h 532: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h 533: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,24,-1,
14'h 534: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,-1,
14'h 535: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,29,-1,
14'h 536: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //25,26,27,28,29,30,31,-1,
14'h 537: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,32,33,-1,
14'h 540: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h 541: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,24,-1,
14'h 542: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h 543: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,27,28,-1,
14'h 544: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //25,26,27,28,29,30,31,-1,
14'h 545: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,32,33,-1,
14'h 546: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //29,30,31,32,33,34,35,-1,
14'h 547: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //31,32,33,34,35,36,37,-1,
14'h 550: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h 551: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,27,28,-1,
14'h 552: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,30,-1,
14'h 553: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //26,27,28,29,30,31,32,-1,
14'h 554: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //29,30,31,32,33,34,35,-1,
14'h 555: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //31,32,33,34,35,36,37,-1,
14'h 556: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //33,34,35,36,37,38,39,-1,
14'h 557: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //35,36,37,38,39,40,41,-1,
14'h 560: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,30,-1,
14'h 561: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //26,27,28,29,30,31,32,-1,
14'h 562: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,34,-1,
14'h 563: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //30,31,32,33,34,35,36,-1,
14'h 564: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //33,34,35,36,37,38,39,-1,
14'h 565: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //35,36,37,38,39,40,41,-1,
14'h 566: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //37,38,39,40,41,42,43,-1,
14'h 567: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //39,40,41,42,43,44,45,-1,
14'h 570: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,34,-1,
14'h 571: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //30,31,32,33,34,35,36,-1,
14'h 572: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //32,33,34,35,36,37,38,-1,
14'h 573: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //34,35,36,37,38,39,40,-1,
14'h 574: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //37,38,39,40,41,42,43,-1,
14'h 575: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //39,40,41,42,43,44,45,-1,
14'h 576: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,-1,
14'h 577: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 3; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 7; adrVal[7]= 7;   end //43,44,45,46,47,48,49,-1,
14'h 600: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,6,-1,
14'h 601: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,7,8,-1,
14'h 602: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,9,-1,
14'h 603: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h 604: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,11,12,-1,
14'h 605: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h 606: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h 607: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h 610: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,10,-1,
14'h 611: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,11,12,-1,
14'h 612: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h 613: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h 614: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h 615: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h 616: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h 617: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h 620: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h 621: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h 622: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h 623: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h 624: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h 625: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h 626: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,24,-1,
14'h 627: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h 630: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h 631: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h 632: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h 633: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h 634: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,24,-1,
14'h 635: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h 636: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,27,28,-1,
14'h 637: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,29,-1,
14'h 640: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h 641: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,24,-1,
14'h 642: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h 643: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,-1,
14'h 644: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,27,28,-1,
14'h 645: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,30,-1,
14'h 646: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //26,27,28,29,30,31,32,-1,
14'h 647: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,32,33,-1,
14'h 650: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h 651: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,27,28,-1,
14'h 652: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,29,-1,
14'h 653: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //25,26,27,28,29,30,31,-1,
14'h 654: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //26,27,28,29,30,31,32,-1,
14'h 655: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,34,-1,
14'h 656: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //30,31,32,33,34,35,36,-1,
14'h 657: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //31,32,33,34,35,36,37,-1,
14'h 660: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,30,-1,
14'h 661: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //26,27,28,29,30,31,32,-1,
14'h 662: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,32,33,-1,
14'h 663: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //29,30,31,32,33,34,35,-1,
14'h 664: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //30,31,32,33,34,35,36,-1,
14'h 665: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //32,33,34,35,36,37,38,-1,
14'h 666: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //34,35,36,37,38,39,40,-1,
14'h 667: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //35,36,37,38,39,40,41,-1,
14'h 670: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,34,-1,
14'h 671: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //30,31,32,33,34,35,36,-1,
14'h 672: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //31,32,33,34,35,36,37,-1,
14'h 673: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //33,34,35,36,37,38,39,-1,
14'h 674: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //34,35,36,37,38,39,40,-1,
14'h 675: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //36,37,38,39,40,41,42,-1,
14'h 676: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //38,39,40,41,42,43,44,-1,
14'h 677: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 3; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 7;   end //39,40,41,42,43,44,45,-1,
14'h 700: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,-1,-1,
14'h 701: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,-1,-1,
14'h 702: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,7,-1,-1,
14'h 703: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,-1,-1,
14'h 704: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,-1,-1,
14'h 705: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h 706: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h 707: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h 710: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,-1,-1,
14'h 711: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h 712: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,11,-1,-1,
14'h 713: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h 714: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h 715: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h 716: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h 717: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h 720: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h 721: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h 722: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,-1,-1,
14'h 723: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h 724: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h 725: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h 726: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h 727: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h 730: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h 731: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h 732: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,-1,-1,
14'h 733: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h 734: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h 735: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h 736: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h 737: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h 740: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h 741: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h 742: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,-1,-1,
14'h 743: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h 744: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h 745: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h 746: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,-1,-1,
14'h 747: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,-1,-1,
14'h 750: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h 751: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h 752: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,27,-1,-1,
14'h 753: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,-1,-1,
14'h 754: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,-1,-1,
14'h 755: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //25,26,27,28,29,30,-1,-1,
14'h 756: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,32,-1,-1,
14'h 757: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,-1,-1,
14'h 760: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,-1,-1,
14'h 761: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //25,26,27,28,29,30,-1,-1,
14'h 762: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //26,27,28,29,30,31,-1,-1,
14'h 763: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,32,-1,-1,
14'h 764: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,-1,-1,
14'h 765: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //29,30,31,32,33,34,-1,-1,
14'h 766: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //31,32,33,34,35,36,-1,-1,
14'h 767: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //32,33,34,35,36,37,-1,-1,
14'h 770: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,-1,-1,
14'h 771: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //29,30,31,32,33,34,-1,-1,
14'h 772: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //30,31,32,33,34,35,-1,-1,
14'h 773: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //31,32,33,34,35,36,-1,-1,
14'h 774: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //32,33,34,35,36,37,-1,-1,
14'h 775: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //33,34,35,36,37,38,-1,-1,
14'h 776: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //35,36,37,38,39,40,-1,-1,
14'h 777: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 3; adrVal[6]= 3; adrVal[7]= 3;   end //36,37,38,39,40,41,-1,-1,
14'h 800: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,-1,-1,
14'h 801: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,-1,-1,
14'h 802: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,-1,-1,
14'h 803: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,7,-1,-1,
14'h 804: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,7,-1,-1,
14'h 805: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,-1,-1,
14'h 806: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,-1,-1,
14'h 807: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,-1,-1,
14'h 810: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,-1,-1,
14'h 811: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,-1,-1,
14'h 812: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h 813: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,11,-1,-1,
14'h 814: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,11,-1,-1,
14'h 815: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h 816: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h 817: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h 820: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h 821: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h 822: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h 823: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,-1,-1,
14'h 824: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,-1,-1,
14'h 825: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h 826: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h 827: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h 830: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h 831: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h 832: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h 833: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,-1,-1,
14'h 834: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,-1,-1,
14'h 835: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h 836: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h 837: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h 840: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h 841: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h 842: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h 843: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,-1,-1,
14'h 844: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,-1,-1,
14'h 845: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h 846: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h 847: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h 850: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h 851: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h 852: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h 853: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,27,-1,-1,
14'h 854: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,27,-1,-1,
14'h 855: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,-1,-1,
14'h 856: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,-1,-1,
14'h 857: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,-1,-1,
14'h 860: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,-1,-1,
14'h 861: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,-1,-1,
14'h 862: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //25,26,27,28,29,30,-1,-1,
14'h 863: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //26,27,28,29,30,31,-1,-1,
14'h 864: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //26,27,28,29,30,31,-1,-1,
14'h 865: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,32,-1,-1,
14'h 866: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,32,-1,-1,
14'h 867: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,-1,-1,
14'h 870: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,-1,-1,
14'h 871: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,-1,-1,
14'h 872: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //29,30,31,32,33,34,-1,-1,
14'h 873: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //30,31,32,33,34,35,-1,-1,
14'h 874: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //30,31,32,33,34,35,-1,-1,
14'h 875: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //31,32,33,34,35,36,-1,-1,
14'h 876: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //31,32,33,34,35,36,-1,-1,
14'h 877: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 3; adrVal[7]= 3;   end //32,33,34,35,36,37,-1,-1,
14'h 900: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,-1,-1,
14'h 901: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,-1,-1,
14'h 902: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,-1,-1,
14'h 903: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,-1,-1,
14'h 904: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,-1,-1,
14'h 905: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,-1,-1,
14'h 906: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,-1,-1,
14'h 907: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,-1,-1,
14'h 910: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,-1,-1,
14'h 911: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,-1,-1,
14'h 912: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,-1,-1,
14'h 913: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,-1,-1,
14'h 914: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h 915: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h 916: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h 917: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h 920: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h 921: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h 922: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h 923: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h 924: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h 925: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h 926: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h 927: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h 930: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h 931: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h 932: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h 933: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h 934: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h 935: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h 936: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h 937: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h 940: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h 941: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h 942: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h 943: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h 944: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h 945: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h 946: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h 947: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h 950: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h 951: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h 952: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h 953: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h 954: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h 955: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h 956: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h 957: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h 960: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,-1,-1,
14'h 961: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,-1,-1,
14'h 962: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,-1,-1,
14'h 963: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,-1,-1,
14'h 964: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //25,26,27,28,29,30,-1,-1,
14'h 965: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //25,26,27,28,29,30,-1,-1,
14'h 966: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //25,26,27,28,29,30,-1,-1,
14'h 967: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //25,26,27,28,29,30,-1,-1,
14'h 970: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,-1,-1,
14'h 971: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,-1,-1,
14'h 972: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,-1,-1,
14'h 973: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,32,33,-1,-1,
14'h 974: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //29,30,31,32,33,34,-1,-1,
14'h 975: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //29,30,31,32,33,34,-1,-1,
14'h 976: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //29,30,31,32,33,34,-1,-1,
14'h 977: begin  adrVal[0]= 1; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //29,30,31,32,33,34,-1,-1,
14'h a00: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,0,1,2,3,
14'h a01: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,6,7,
14'h a02: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,8,9,10,11,
14'h a03: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,12,13,14,15,
14'h a04: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,-1,-1,-1,-1,
14'h a05: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,-1,-1,-1,-1,
14'h a06: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,-1,-1,-1,-1,
14'h a07: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,-1,-1,-1,-1,
14'h a10: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,-1,-1,-1,-1,
14'h a11: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,-1,-1,-1,-1,
14'h a12: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,-1,-1,-1,-1,
14'h a13: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,-1,-1,-1,-1,
14'h a14: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,-1,-1,-1,-1,
14'h a15: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,-1,-1,-1,-1,
14'h a16: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,-1,-1,-1,-1,
14'h a17: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,-1,-1,-1,-1,
14'h a20: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h a21: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h a22: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h a23: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h a24: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h a25: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h a26: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h a27: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h a30: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h a31: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h a32: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h a33: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h a34: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h a35: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h a36: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h a37: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h a40: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h a41: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h a42: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h a43: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h a44: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h a45: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h a46: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h a47: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h a50: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h a51: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h a52: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h a53: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h a54: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h a55: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h a56: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h a57: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h a60: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,-1,-1,-1,-1,
14'h a61: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,-1,-1,-1,-1,
14'h a62: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,-1,-1,-1,-1,
14'h a63: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,-1,-1,-1,-1,
14'h a64: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,-1,-1,-1,-1,
14'h a65: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,-1,-1,-1,-1,
14'h a66: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,-1,-1,-1,-1,
14'h a67: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,-1,-1,-1,-1,
14'h a70: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,-1,-1,-1,-1,
14'h a71: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,-1,-1,-1,-1,
14'h a72: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,-1,-1,-1,-1,
14'h a73: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,-1,-1,-1,-1,
14'h a74: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,-1,-1,-1,-1,
14'h a75: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,-1,-1,-1,-1,
14'h a76: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,-1,-1,-1,-1,
14'h a77: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //28,29,30,31,-1,-1,-1,-1,
14'h b00: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,-1,-1,-1,
14'h b01: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,-1,-1,-1,
14'h b02: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,-1,-1,-1,
14'h b03: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,-1,-1,-1,
14'h b04: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //15,99,0,1,2,-1,-1,-1,
14'h b05: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //15,99,0,1,2,-1,-1,-1,
14'h b06: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //15,99,0,1,2,-1,-1,-1,
14'h b07: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //15,99,0,1,2,-1,-1,-1,
14'h b10: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,-1,-1,-1,
14'h b11: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,-1,-1,-1,
14'h b12: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,-1,-1,-1,
14'h b13: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,-1,-1,-1,
14'h b14: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,-1,-1,-1,
14'h b15: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,-1,-1,-1,
14'h b16: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,-1,-1,-1,
14'h b17: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,-1,-1,-1,
14'h b20: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,-1,-1,-1,
14'h b21: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,-1,-1,-1,
14'h b22: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,-1,-1,-1,
14'h b23: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,-1,-1,-1,
14'h b24: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,-1,-1,-1,
14'h b25: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,-1,-1,-1,
14'h b26: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,-1,-1,-1,
14'h b27: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,-1,-1,-1,
14'h b30: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,-1,-1,-1,
14'h b31: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,-1,-1,-1,
14'h b32: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,-1,-1,-1,
14'h b33: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,-1,-1,-1,
14'h b34: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,-1,-1,-1,
14'h b35: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,-1,-1,-1,
14'h b36: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,-1,-1,-1,
14'h b37: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,-1,-1,-1,
14'h b40: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,-1,-1,-1,
14'h b41: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,-1,-1,-1,
14'h b42: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,-1,-1,-1,
14'h b43: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,-1,-1,-1,
14'h b44: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,-1,-1,-1,
14'h b45: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,-1,-1,-1,
14'h b46: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,-1,-1,-1,
14'h b47: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,-1,-1,-1,
14'h b50: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,-1,-1,-1,
14'h b51: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,-1,-1,-1,
14'h b52: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,-1,-1,-1,
14'h b53: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,-1,-1,-1,
14'h b54: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,-1,-1,-1,
14'h b55: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,-1,-1,-1,
14'h b56: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,-1,-1,-1,
14'h b57: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,-1,-1,-1,
14'h b60: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,-1,-1,-1,
14'h b61: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,-1,-1,-1,
14'h b62: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,-1,-1,-1,
14'h b63: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,-1,-1,-1,
14'h b64: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,-1,-1,-1,
14'h b65: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,-1,-1,-1,
14'h b66: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,-1,-1,-1,
14'h b67: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,-1,-1,-1,
14'h b70: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,-1,-1,-1,
14'h b71: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,-1,-1,-1,
14'h b72: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,-1,-1,-1,
14'h b73: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,-1,-1,-1,
14'h b74: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //26,27,28,29,30,-1,-1,-1,
14'h b75: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //26,27,28,29,30,-1,-1,-1,
14'h b76: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //26,27,28,29,30,-1,-1,-1,
14'h b77: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //26,27,28,29,30,-1,-1,-1,
14'h c00: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,4,-1,-1,
14'h c01: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //5,99,0,1,2,3,-1,-1,
14'h c02: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //5,99,0,1,2,3,-1,-1,
14'h c03: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //12,5,99,0,1,2,-1,-1,
14'h c04: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //18,12,5,99,0,1,-1,-1,
14'h c05: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //18,12,5,99,0,1,-1,-1,
14'h c06: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 1;   end //25,18,12,5,99,0,-1,-1,
14'h c07: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 1;   end //25,18,12,5,99,0,-1,-1,
14'h c10: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,-1,-1,
14'h c11: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,7,-1,-1,
14'h c12: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,7,-1,-1,
14'h c13: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,-1,-1,
14'h c14: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,-1,-1,
14'h c15: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,-1,-1,
14'h c16: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,4,-1,-1,
14'h c17: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,4,-1,-1,
14'h c20: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h c21: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,11,-1,-1,
14'h c22: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,11,-1,-1,
14'h c23: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h c24: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,-1,-1,
14'h c25: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,-1,-1,
14'h c26: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,-1,-1,
14'h c27: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,-1,-1,
14'h c30: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h c31: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,-1,-1,
14'h c32: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,-1,-1,
14'h c33: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h c34: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h c35: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h c36: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h c37: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h c40: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h c41: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,-1,-1,
14'h c42: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,-1,-1,
14'h c43: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h c44: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h c45: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h c46: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h c47: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h c50: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h c51: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,-1,-1,
14'h c52: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,-1,-1,
14'h c53: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h c54: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h c55: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h c56: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h c57: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h c60: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,-1,-1,
14'h c61: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,27,-1,-1,
14'h c62: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,27,-1,-1,
14'h c63: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h c64: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h c65: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h c66: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h c67: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h c70: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //27,28,29,30,31,32,-1,-1,
14'h c71: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //26,27,28,29,30,31,-1,-1,
14'h c72: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //26,27,28,29,30,31,-1,-1,
14'h c73: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //25,26,27,28,29,30,-1,-1,
14'h c74: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,-1,-1,
14'h c75: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,-1,-1,
14'h c76: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,-1,-1,
14'h c77: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,-1,-1,
14'h d00: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //3,99,0,1,2,3,-1,-1,
14'h d01: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //6,3,99,0,1,2,-1,-1,
14'h d02: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //10,6,3,99,0,1,-1,-1,
14'h d03: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //13,10,6,3,99,0,-1,-1,
14'h d04: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //17,13,10,6,3,99,-1,-1,
14'h d05: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //20,17,13,10,6,3,-1,-1,
14'h d06: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //24,20,17,13,10,6,-1,-1,
14'h d07: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //27,24,20,17,13,10,-1,-1,
14'h d10: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,7,-1,-1,
14'h d11: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,-1,-1,
14'h d12: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,-1,-1,
14'h d13: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,4,-1,-1,
14'h d14: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //3,99,0,1,2,3,-1,-1,
14'h d15: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //6,3,99,0,1,2,-1,-1,
14'h d16: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //10,6,3,99,0,1,-1,-1,
14'h d17: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //13,10,6,3,99,0,-1,-1,
14'h d20: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,11,-1,-1,
14'h d21: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h d22: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,-1,-1,
14'h d23: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,-1,-1,
14'h d24: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,7,-1,-1,
14'h d25: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,-1,-1,
14'h d26: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,-1,-1,
14'h d27: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,4,-1,-1,
14'h d30: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,-1,-1,
14'h d31: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h d32: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h d33: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h d34: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,11,-1,-1,
14'h d35: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h d36: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,-1,-1,
14'h d37: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,-1,-1,
14'h d40: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,-1,-1,
14'h d41: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h d42: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h d43: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h d44: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,-1,-1,
14'h d45: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h d46: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h d47: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h d50: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,-1,-1,
14'h d51: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h d52: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h d53: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h d54: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,-1,-1,
14'h d55: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h d56: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h d57: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h d60: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,27,-1,-1,
14'h d61: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h d62: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h d63: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h d64: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,-1,-1,
14'h d65: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h d66: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h d67: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h d70: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //26,27,28,29,30,31,-1,-1,
14'h d71: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //25,26,27,28,29,30,-1,-1,
14'h d72: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,-1,-1,
14'h d73: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,-1,-1,
14'h d74: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,27,-1,-1,
14'h d75: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h d76: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h d77: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h e00: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //1,99,0,1,2,3,4,-1,
14'h e01: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //6,4,1,99,0,1,2,-1,
14'h e02: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //9,6,4,1,99,0,1,-1,
14'h e03: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //14,11,9,6,4,1,99,-1,
14'h e04: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //19,16,14,11,9,6,4,-1,
14'h e05: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //21,19,16,14,11,9,6,-1,
14'h e06: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //26,24,21,19,16,14,11,-1,
14'h e07: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //29,26,24,21,19,16,14,-1,
14'h e10: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,7,8,-1,
14'h e11: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,6,-1,
14'h e12: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,4,5,-1,
14'h e13: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //4,1,99,0,1,2,3,-1,
14'h e14: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //9,6,4,1,99,0,1,-1,
14'h e15: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //11,9,6,4,1,99,0,-1,
14'h e16: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,14,11,9,6,4,1,-1,
14'h e17: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //19,16,14,11,9,6,4,-1,
14'h e20: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,11,12,-1,
14'h e21: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,10,-1,
14'h e22: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,9,-1,
14'h e23: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,7,-1,
14'h e24: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,4,5,-1,
14'h e25: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //1,99,0,1,2,3,4,-1,
14'h e26: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //6,4,1,99,0,1,2,-1,
14'h e27: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //9,6,4,1,99,0,1,-1,
14'h e30: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h e31: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h e32: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h e33: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h e34: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,9,-1,
14'h e35: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,7,8,-1,
14'h e36: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,6,-1,
14'h e37: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,4,5,-1,
14'h e40: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h e41: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h e42: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h e43: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h e44: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h e45: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,11,12,-1,
14'h e46: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,10,-1,
14'h e47: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,9,-1,
14'h e50: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,24,-1,
14'h e51: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h e52: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h e53: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h e54: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h e55: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h e56: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h e57: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h e60: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,27,28,-1,
14'h e61: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h e62: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h e63: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h e64: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h e65: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h e66: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h e67: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h e70: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //26,27,28,29,30,31,32,-1,
14'h e71: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //24,25,26,27,28,29,30,-1,
14'h e72: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,29,-1,
14'h e73: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,-1,
14'h e74: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h e75: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,24,-1,
14'h e76: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h e77: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h f00: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //3,1,99,0,1,2,3,-1,
14'h f01: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //7,5,3,1,99,0,1,-1,
14'h f02: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //10,8,7,5,3,1,99,-1,
14'h f03: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,12,10,8,7,5,3,-1,
14'h f04: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,16,14,12,10,8,7,-1,
14'h f05: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //22,20,18,16,14,12,10,-1,
14'h f06: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //25,23,22,20,18,16,14,-1,
14'h f07: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //29,27,25,23,22,20,18,-1,
14'h f10: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,7,-1,
14'h f11: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,4,5,-1,
14'h f12: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //3,1,99,0,1,2,3,-1,
14'h f13: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //7,5,3,1,99,0,1,-1,
14'h f14: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //10,8,7,5,3,1,99,-1,
14'h f15: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,12,10,8,7,5,3,-1,
14'h f16: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,16,14,12,10,8,7,-1,
14'h f17: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //22,20,18,16,14,12,10,-1,
14'h f20: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h f21: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,9,-1,
14'h f22: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,7,-1,
14'h f23: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,4,5,-1,
14'h f24: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //3,1,99,0,1,2,3,-1,
14'h f25: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //7,5,3,1,99,0,1,-1,
14'h f26: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //10,8,7,5,3,1,99,-1,
14'h f27: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,12,10,8,7,5,3,-1,
14'h f30: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h f31: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h f32: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h f33: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,9,-1,
14'h f34: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,7,-1,
14'h f35: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,4,5,-1,
14'h f36: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //3,1,99,0,1,2,3,-1,
14'h f37: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //7,5,3,1,99,0,1,-1,
14'h f40: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h f41: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h f42: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h f43: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h f44: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h f45: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,9,-1,
14'h f46: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,7,-1,
14'h f47: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,4,5,-1,
14'h f50: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h f51: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h f52: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h f53: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h f54: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h f55: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h f56: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h f57: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,9,-1,
14'h f60: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,-1,
14'h f61: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h f62: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h f63: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h f64: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h f65: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h f66: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h f67: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h f70: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //25,26,27,28,29,30,31,-1,
14'h f71: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,24,25,26,27,28,29,-1,
14'h f72: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,-1,
14'h f73: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h f74: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h f75: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h f76: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h f77: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h1000: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //2,1,99,0,1,2,3,-1,
14'h1001: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //7,5,4,2,1,99,0,-1,
14'h1002: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,8,7,5,4,2,1,-1,
14'h1003: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,13,11,10,8,7,5,-1,
14'h1004: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //19,17,16,14,13,11,10,-1,
14'h1005: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //22,20,19,17,16,14,13,-1,
14'h1006: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //26,25,23,22,20,19,17,-1,
14'h1007: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //29,28,26,25,23,22,20,-1,
14'h1010: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,7,-1,
14'h1011: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //1,99,0,1,2,3,4,-1,
14'h1012: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //4,2,1,99,0,1,2,-1,
14'h1013: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //8,7,5,4,2,1,99,-1,
14'h1014: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,11,10,8,7,5,4,-1,
14'h1015: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,14,13,11,10,8,7,-1,
14'h1016: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //20,19,17,16,14,13,11,-1,
14'h1017: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //23,22,20,19,17,16,14,-1,
14'h1020: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h1021: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,7,8,-1,
14'h1022: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,6,-1,
14'h1023: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //2,1,99,0,1,2,3,-1,
14'h1024: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //7,5,4,2,1,99,0,-1,
14'h1025: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,8,7,5,4,2,1,-1,
14'h1026: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,13,11,10,8,7,5,-1,
14'h1027: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,16,14,13,11,10,8,-1,
14'h1030: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h1031: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,11,12,-1,
14'h1032: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,10,-1,
14'h1033: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,7,-1,
14'h1034: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //1,99,0,1,2,3,4,-1,
14'h1035: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //4,2,1,99,0,1,2,-1,
14'h1036: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //8,7,5,4,2,1,99,-1,
14'h1037: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,10,8,7,5,4,2,-1,
14'h1040: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h1041: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h1042: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h1043: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h1044: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,7,8,-1,
14'h1045: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,6,-1,
14'h1046: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //2,1,99,0,1,2,3,-1,
14'h1047: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //5,4,2,1,99,0,1,-1,
14'h1050: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h1051: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h1052: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h1053: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h1054: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,11,12,-1,
14'h1055: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,10,-1,
14'h1056: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,7,-1,
14'h1057: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,4,5,-1,
14'h1060: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,-1,
14'h1061: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,24,-1,
14'h1062: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h1063: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h1064: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h1065: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h1066: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h1067: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,9,-1,
14'h1070: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //25,26,27,28,29,30,31,-1,
14'h1071: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,23,24,25,26,27,28,-1,
14'h1072: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h1073: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h1074: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h1075: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h1076: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h1077: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h1100: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //3,1,0,99,0,1,2,3,
14'h1101: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //6,5,4,3,1,0,99,0,
14'h1102: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,9,8,6,5,4,3,1,
14'h1103: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,13,11,10,9,8,6,5,
14'h1104: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //19,17,16,15,14,13,11,10,
14'h1105: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //22,21,20,19,17,16,15,14,
14'h1106: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //26,25,24,22,21,20,19,17,
14'h1107: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //30,29,27,26,25,24,22,21,
14'h1110: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,6,7,
14'h1111: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //1,0,99,0,1,2,3,4,
14'h1112: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //5,4,3,1,0,99,0,1,
14'h1113: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,8,6,5,4,3,1,0,
14'h1114: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,13,11,10,9,8,6,5,
14'h1115: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,16,15,14,13,11,10,9,
14'h1116: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //21,20,19,17,16,15,14,13,
14'h1117: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //25,24,22,21,20,19,17,16,
14'h1120: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,10,11,
14'h1121: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,7,8,
14'h1122: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,99,0,1,2,3,4,5,
14'h1123: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //4,3,1,0,99,0,1,2,
14'h1124: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,8,6,5,4,3,1,0,
14'h1125: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,11,10,9,8,6,5,4,
14'h1126: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,15,14,13,11,10,9,8,
14'h1127: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //20,19,17,16,15,14,13,11,
14'h1130: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,14,15,
14'h1131: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,11,12,
14'h1132: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,7,8,9,
14'h1133: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,4,5,6,
14'h1134: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //4,3,1,0,99,0,1,2,
14'h1135: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //8,6,5,4,3,1,0,99,
14'h1136: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,10,9,8,6,5,4,3,
14'h1137: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,14,13,11,10,9,8,6,
14'h1140: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,19,
14'h1141: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,16,
14'h1142: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //6,7,8,9,10,11,12,13,
14'h1143: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,9,10,
14'h1144: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //99,0,1,2,3,4,5,6,
14'h1145: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //3,1,0,99,0,1,2,3,
14'h1146: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //6,5,4,3,1,0,99,0,
14'h1147: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,9,8,6,5,4,3,1,
14'h1150: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,23,
14'h1151: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,20,
14'h1152: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,17,
14'h1153: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,13,14,
14'h1154: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //3,4,5,6,7,8,9,10,
14'h1155: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,6,7,
14'h1156: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //1,0,99,0,1,2,3,4,
14'h1157: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //5,4,3,1,0,99,0,1,
14'h1160: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //20,21,22,23,24,25,26,27,
14'h1161: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,23,24,
14'h1162: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,21,
14'h1163: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,18,
14'h1164: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //7,8,9,10,11,12,13,14,
14'h1165: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //4,5,6,7,8,9,10,11,
14'h1166: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //1,2,3,4,5,6,7,8,
14'h1167: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,99,0,1,2,3,4,5,
14'h1170: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 3;   end //24,25,26,27,28,29,30,31,
14'h1171: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,22,23,24,25,26,27,28,
14'h1172: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,23,24,25,
14'h1173: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,22,
14'h1174: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,18,
14'h1175: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //8,9,10,11,12,13,14,15,
14'h1176: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //5,6,7,8,9,10,11,12,
14'h1177: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //2,3,4,5,6,7,8,9,
14'h1200: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //2,1,0,99,0,1,2,3,
14'h1201: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //6,5,4,3,2,1,0,99,
14'h1202: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //10,9,8,7,6,5,4,3,
14'h1203: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //14,13,12,11,10,9,8,7,
14'h1204: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //18,17,16,15,14,13,12,11,
14'h1205: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,21,20,19,18,17,16,15,
14'h1206: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //26,25,24,23,22,21,20,19,
14'h1207: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //30,29,28,27,26,25,24,23,
14'h1210: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,7,
14'h1211: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //2,1,0,99,0,1,2,3,
14'h1212: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //6,5,4,3,2,1,0,99,
14'h1213: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //10,9,8,7,6,5,4,3,
14'h1214: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //14,13,12,11,10,9,8,7,
14'h1215: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //18,17,16,15,14,13,12,11,
14'h1216: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,21,20,19,18,17,16,15,
14'h1217: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //26,25,24,23,22,21,20,19,
14'h1220: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,11,
14'h1221: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,7,
14'h1222: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //2,1,0,99,0,1,2,3,
14'h1223: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //6,5,4,3,2,1,0,99,
14'h1224: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //10,9,8,7,6,5,4,3,
14'h1225: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //14,13,12,11,10,9,8,7,
14'h1226: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //18,17,16,15,14,13,12,11,
14'h1227: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,21,20,19,18,17,16,15,
14'h1230: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,15,
14'h1231: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,11,
14'h1232: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,7,
14'h1233: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //2,1,0,99,0,1,2,3,
14'h1234: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //6,5,4,3,2,1,0,99,
14'h1235: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //10,9,8,7,6,5,4,3,
14'h1236: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //14,13,12,11,10,9,8,7,
14'h1237: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //18,17,16,15,14,13,12,11,
14'h1240: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,19,
14'h1241: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,15,
14'h1242: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,11,
14'h1243: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,7,
14'h1244: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //2,1,0,99,0,1,2,3,
14'h1245: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //6,5,4,3,2,1,0,99,
14'h1246: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //10,9,8,7,6,5,4,3,
14'h1247: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //14,13,12,11,10,9,8,7,
14'h1250: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //16,17,18,19,20,21,22,23,
14'h1251: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,19,
14'h1252: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,15,
14'h1253: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,11,
14'h1254: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,7,
14'h1255: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //2,1,0,99,0,1,2,3,
14'h1256: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //6,5,4,3,2,1,0,99,
14'h1257: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //10,9,8,7,6,5,4,3,
14'h1260: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //20,21,22,23,24,25,26,27,
14'h1261: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //16,17,18,19,20,21,22,23,
14'h1262: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,19,
14'h1263: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,15,
14'h1264: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,11,
14'h1265: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,7,
14'h1266: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //2,1,0,99,0,1,2,3,
14'h1267: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //6,5,4,3,2,1,0,99,
14'h1270: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,30,31,
14'h1271: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //20,21,22,23,24,25,26,27,
14'h1272: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //16,17,18,19,20,21,22,23,
14'h1273: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,19,
14'h1274: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,15,
14'h1275: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,11,
14'h1276: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,7,
14'h1277: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //2,1,0,99,0,1,2,3,
14'h1300: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //3,1,0,99,0,1,2,3,
14'h1301: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //6,5,4,3,1,0,99,0,
14'h1302: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //10,9,8,6,5,4,3,1,
14'h1303: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //14,13,11,10,9,8,6,5,
14'h1304: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //19,17,16,15,14,13,11,10,
14'h1305: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,21,20,19,17,16,15,14,
14'h1306: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //26,25,24,22,21,20,19,17,
14'h1307: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //30,29,27,26,25,24,22,21,
14'h1310: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,7,
14'h1311: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //1,0,99,0,1,2,3,4,
14'h1312: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //5,4,3,1,0,99,0,1,
14'h1313: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //9,8,6,5,4,3,1,0,
14'h1314: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //14,13,11,10,9,8,6,5,
14'h1315: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //17,16,15,14,13,11,10,9,
14'h1316: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //21,20,19,17,16,15,14,13,
14'h1317: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //25,24,22,21,20,19,17,16,
14'h1320: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,11,
14'h1321: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,7,8,
14'h1322: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //0,99,0,1,2,3,4,5,
14'h1323: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //4,3,1,0,99,0,1,2,
14'h1324: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //9,8,6,5,4,3,1,0,
14'h1325: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //13,11,10,9,8,6,5,4,
14'h1326: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //16,15,14,13,11,10,9,8,
14'h1327: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //20,19,17,16,15,14,13,11,
14'h1330: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,15,
14'h1331: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,11,12,
14'h1332: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,7,8,9,
14'h1333: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,4,5,6,
14'h1334: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //4,3,1,0,99,0,1,2,
14'h1335: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //8,6,5,4,3,1,0,99,
14'h1336: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //11,10,9,8,6,5,4,3,
14'h1337: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //15,14,13,11,10,9,8,6,
14'h1340: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,19,
14'h1341: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,16,
14'h1342: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,11,12,13,
14'h1343: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,9,10,
14'h1344: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,4,5,6,
14'h1345: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //3,1,0,99,0,1,2,3,
14'h1346: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //6,5,4,3,1,0,99,0,
14'h1347: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //10,9,8,6,5,4,3,1,
14'h1350: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //16,17,18,19,20,21,22,23,
14'h1351: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,20,
14'h1352: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,17,
14'h1353: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,13,14,
14'h1354: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,9,10,
14'h1355: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,7,
14'h1356: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //1,0,99,0,1,2,3,4,
14'h1357: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //5,4,3,1,0,99,0,1,
14'h1360: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //20,21,22,23,24,25,26,27,
14'h1361: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,24,
14'h1362: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,21,
14'h1363: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,18,
14'h1364: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,13,14,
14'h1365: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,11,
14'h1366: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,7,8,
14'h1367: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //0,99,0,1,2,3,4,5,
14'h1370: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,30,31,
14'h1371: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,28,
14'h1372: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,24,25,
14'h1373: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,22,
14'h1374: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,18,
14'h1375: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,15,
14'h1376: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,11,12,
14'h1377: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,7,8,9,
14'h1400: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //2,1,99,0,1,2,3,-1,
14'h1401: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //7,5,4,2,1,99,0,-1,
14'h1402: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //10,8,7,5,4,2,1,-1,
14'h1403: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //14,13,11,10,8,7,5,-1,
14'h1404: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //19,17,16,14,13,11,10,-1,
14'h1405: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //22,20,19,17,16,14,13,-1,
14'h1406: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //26,25,23,22,20,19,17,-1,
14'h1407: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //29,28,26,25,23,22,20,-1,
14'h1410: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,7,-1,
14'h1411: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //1,99,0,1,2,3,4,-1,
14'h1412: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //4,2,1,99,0,1,2,-1,
14'h1413: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //8,7,5,4,2,1,99,-1,
14'h1414: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //13,11,10,8,7,5,4,-1,
14'h1415: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //16,14,13,11,10,8,7,-1,
14'h1416: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //20,19,17,16,14,13,11,-1,
14'h1417: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //23,22,20,19,17,16,14,-1,
14'h1420: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h1421: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,7,8,-1,
14'h1422: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,-1,
14'h1423: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //2,1,99,0,1,2,3,-1,
14'h1424: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //7,5,4,2,1,99,0,-1,
14'h1425: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //10,8,7,5,4,2,1,-1,
14'h1426: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //14,13,11,10,8,7,5,-1,
14'h1427: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //17,16,14,13,11,10,8,-1,
14'h1430: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h1431: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,11,12,-1,
14'h1432: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,-1,
14'h1433: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,7,-1,
14'h1434: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //1,99,0,1,2,3,4,-1,
14'h1435: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //4,2,1,99,0,1,2,-1,
14'h1436: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //8,7,5,4,2,1,99,-1,
14'h1437: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //11,10,8,7,5,4,2,-1,
14'h1440: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h1441: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h1442: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h1443: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h1444: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,7,8,-1,
14'h1445: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,-1,
14'h1446: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //2,1,99,0,1,2,3,-1,
14'h1447: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //5,4,2,1,99,0,1,-1,
14'h1450: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h1451: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h1452: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h1453: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h1454: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,11,12,-1,
14'h1455: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,-1,
14'h1456: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,7,-1,
14'h1457: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,4,5,-1,
14'h1460: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,-1,
14'h1461: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,24,-1,
14'h1462: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h1463: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h1464: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h1465: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h1466: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h1467: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,9,-1,
14'h1470: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,31,-1,
14'h1471: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //22,23,24,25,26,27,28,-1,
14'h1472: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h1473: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h1474: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h1475: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h1476: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h1477: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h1500: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //3,1,99,0,1,2,3,-1,
14'h1501: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //7,5,3,1,99,0,1,-1,
14'h1502: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //10,8,7,5,3,1,99,-1,
14'h1503: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //14,12,10,8,7,5,3,-1,
14'h1504: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //18,16,14,12,10,8,7,-1,
14'h1505: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //22,20,18,16,14,12,10,-1,
14'h1506: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //25,23,22,20,18,16,14,-1,
14'h1507: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //29,27,25,23,22,20,18,-1,
14'h1510: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,7,-1,
14'h1511: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,4,5,-1,
14'h1512: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //3,1,99,0,1,2,3,-1,
14'h1513: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //7,5,3,1,99,0,1,-1,
14'h1514: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //10,8,7,5,3,1,99,-1,
14'h1515: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //14,12,10,8,7,5,3,-1,
14'h1516: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //18,16,14,12,10,8,7,-1,
14'h1517: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //22,20,18,16,14,12,10,-1,
14'h1520: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h1521: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,9,-1,
14'h1522: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,7,-1,
14'h1523: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,4,5,-1,
14'h1524: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //3,1,99,0,1,2,3,-1,
14'h1525: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //7,5,3,1,99,0,1,-1,
14'h1526: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //10,8,7,5,3,1,99,-1,
14'h1527: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //14,12,10,8,7,5,3,-1,
14'h1530: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h1531: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h1532: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h1533: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,9,-1,
14'h1534: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,7,-1,
14'h1535: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,4,5,-1,
14'h1536: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //3,1,99,0,1,2,3,-1,
14'h1537: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //7,5,3,1,99,0,1,-1,
14'h1540: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h1541: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h1542: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h1543: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h1544: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h1545: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,9,-1,
14'h1546: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,7,-1,
14'h1547: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,4,5,-1,
14'h1550: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h1551: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h1552: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h1553: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h1554: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h1555: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h1556: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h1557: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,9,-1,
14'h1560: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,-1,
14'h1561: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h1562: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h1563: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h1564: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h1565: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h1566: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h1567: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h1570: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,31,-1,
14'h1571: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,29,-1,
14'h1572: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,-1,
14'h1573: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h1574: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h1575: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h1576: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h1577: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h1600: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //1,99,0,1,2,3,4,-1,
14'h1601: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //6,4,1,99,0,1,2,-1,
14'h1602: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //9,6,4,1,99,0,1,-1,
14'h1603: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //14,11,9,6,4,1,99,-1,
14'h1604: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //19,16,14,11,9,6,4,-1,
14'h1605: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //21,19,16,14,11,9,6,-1,
14'h1606: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //26,24,21,19,16,14,11,-1,
14'h1607: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //29,26,24,21,19,16,14,-1,
14'h1610: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,7,8,-1,
14'h1611: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,-1,
14'h1612: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,4,5,-1,
14'h1613: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //4,1,99,0,1,2,3,-1,
14'h1614: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //9,6,4,1,99,0,1,-1,
14'h1615: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //11,9,6,4,1,99,0,-1,
14'h1616: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //16,14,11,9,6,4,1,-1,
14'h1617: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //19,16,14,11,9,6,4,-1,
14'h1620: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,11,12,-1,
14'h1621: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,-1,
14'h1622: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,9,-1,
14'h1623: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,7,-1,
14'h1624: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,4,5,-1,
14'h1625: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //1,99,0,1,2,3,4,-1,
14'h1626: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //6,4,1,99,0,1,2,-1,
14'h1627: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //9,6,4,1,99,0,1,-1,
14'h1630: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h1631: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h1632: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h1633: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h1634: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,9,-1,
14'h1635: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,7,8,-1,
14'h1636: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,-1,
14'h1637: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,4,5,-1,
14'h1640: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h1641: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h1642: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h1643: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h1644: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h1645: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,11,12,-1,
14'h1646: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,-1,
14'h1647: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,9,-1,
14'h1650: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,24,-1,
14'h1651: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h1652: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h1653: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h1654: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h1655: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h1656: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h1657: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h1660: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //22,23,24,25,26,27,28,-1,
14'h1661: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h1662: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h1663: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h1664: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h1665: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h1666: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h1667: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h1670: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,31,32,-1,
14'h1671: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,30,-1,
14'h1672: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,29,-1,
14'h1673: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,-1,
14'h1674: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h1675: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,24,-1,
14'h1676: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h1677: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h1700: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //3,99,0,1,2,3,-1,-1,
14'h1701: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //6,3,99,0,1,2,-1,-1,
14'h1702: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //10,6,3,99,0,1,-1,-1,
14'h1703: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //13,10,6,3,99,0,-1,-1,
14'h1704: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //17,13,10,6,3,99,-1,-1,
14'h1705: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //20,17,13,10,6,3,-1,-1,
14'h1706: begin  adrVal[0]= 7; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //24,20,17,13,10,6,-1,-1,
14'h1707: begin  adrVal[0]= 1; adrVal[1]= 1; adrVal[2]= 1; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //27,24,20,17,13,10,-1,-1,
14'h1710: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,7,-1,-1,
14'h1711: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,-1,-1,
14'h1712: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,-1,-1,
14'h1713: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,4,-1,-1,
14'h1714: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //3,99,0,1,2,3,-1,-1,
14'h1715: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //6,3,99,0,1,2,-1,-1,
14'h1716: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //10,6,3,99,0,1,-1,-1,
14'h1717: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //13,10,6,3,99,0,-1,-1,
14'h1720: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,11,-1,-1,
14'h1721: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h1722: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,-1,-1,
14'h1723: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,-1,-1,
14'h1724: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,7,-1,-1,
14'h1725: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,-1,-1,
14'h1726: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,-1,-1,
14'h1727: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,4,-1,-1,
14'h1730: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,-1,-1,
14'h1731: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h1732: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h1733: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h1734: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,11,-1,-1,
14'h1735: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h1736: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,-1,-1,
14'h1737: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,-1,-1,
14'h1740: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,-1,-1,
14'h1741: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h1742: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h1743: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h1744: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,-1,-1,
14'h1745: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h1746: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h1747: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h1750: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,-1,-1,
14'h1751: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h1752: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h1753: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h1754: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,-1,-1,
14'h1755: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h1756: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h1757: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h1760: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //22,23,24,25,26,27,-1,-1,
14'h1761: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h1762: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h1763: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h1764: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,-1,-1,
14'h1765: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h1766: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h1767: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h1770: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,31,-1,-1,
14'h1771: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,-1,-1,
14'h1772: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,-1,-1,
14'h1773: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,-1,-1,
14'h1774: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //22,23,24,25,26,27,-1,-1,
14'h1775: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h1776: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h1777: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h1800: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,4,-1,-1,
14'h1801: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //5,99,0,1,2,3,-1,-1,
14'h1802: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //5,99,0,1,2,3,-1,-1,
14'h1803: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //12,5,99,0,1,2,-1,-1,
14'h1804: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //18,12,5,99,0,1,-1,-1,
14'h1805: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //18,12,5,99,0,1,-1,-1,
14'h1806: begin  adrVal[0]= 0; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //25,18,12,5,99,0,-1,-1,
14'h1807: begin  adrVal[0]= 0; adrVal[1]= 1; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //25,18,12,5,99,0,-1,-1,
14'h1810: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,-1,-1,
14'h1811: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,7,-1,-1,
14'h1812: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,7,-1,-1,
14'h1813: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,-1,-1,
14'h1814: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,-1,-1,
14'h1815: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,-1,-1,
14'h1816: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,4,-1,-1,
14'h1817: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,4,-1,-1,
14'h1820: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h1821: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,11,-1,-1,
14'h1822: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,11,-1,-1,
14'h1823: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h1824: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,-1,-1,
14'h1825: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,-1,-1,
14'h1826: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,-1,-1,
14'h1827: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,-1,-1,
14'h1830: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h1831: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,-1,-1,
14'h1832: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,-1,-1,
14'h1833: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h1834: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h1835: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h1836: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h1837: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h1840: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h1841: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,-1,-1,
14'h1842: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,-1,-1,
14'h1843: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h1844: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h1845: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h1846: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h1847: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h1850: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h1851: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,-1,-1,
14'h1852: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,-1,-1,
14'h1853: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h1854: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h1855: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h1856: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h1857: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h1860: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,-1,-1,
14'h1861: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //22,23,24,25,26,27,-1,-1,
14'h1862: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //22,23,24,25,26,27,-1,-1,
14'h1863: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h1864: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h1865: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h1866: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h1867: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h1870: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,32,-1,-1,
14'h1871: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,31,-1,-1,
14'h1872: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,31,-1,-1,
14'h1873: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,-1,-1,
14'h1874: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,-1,-1,
14'h1875: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,-1,-1,
14'h1876: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,-1,-1,
14'h1877: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,-1,-1,
14'h1900: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,-1,-1,-1,
14'h1901: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,-1,-1,-1,
14'h1902: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,-1,-1,-1,
14'h1903: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //99,0,1,2,3,-1,-1,-1,
14'h1904: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //15,99,0,1,2,-1,-1,-1,
14'h1905: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //15,99,0,1,2,-1,-1,-1,
14'h1906: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //15,99,0,1,2,-1,-1,-1,
14'h1907: begin  adrVal[0]= 0; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 1;   end //15,99,0,1,2,-1,-1,-1,
14'h1910: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,-1,-1,-1,
14'h1911: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,-1,-1,-1,
14'h1912: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,-1,-1,-1,
14'h1913: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,-1,-1,-1,
14'h1914: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,-1,-1,-1,
14'h1915: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,-1,-1,-1,
14'h1916: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,-1,-1,-1,
14'h1917: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,-1,-1,-1,
14'h1920: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,-1,-1,-1,
14'h1921: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,-1,-1,-1,
14'h1922: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,-1,-1,-1,
14'h1923: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,-1,-1,-1,
14'h1924: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,-1,-1,-1,
14'h1925: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,-1,-1,-1,
14'h1926: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,-1,-1,-1,
14'h1927: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,-1,-1,-1,
14'h1930: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,-1,-1,-1,
14'h1931: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,-1,-1,-1,
14'h1932: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,-1,-1,-1,
14'h1933: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,-1,-1,-1,
14'h1934: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,-1,-1,-1,
14'h1935: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,-1,-1,-1,
14'h1936: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,-1,-1,-1,
14'h1937: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,-1,-1,-1,
14'h1940: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,-1,-1,-1,
14'h1941: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,-1,-1,-1,
14'h1942: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,-1,-1,-1,
14'h1943: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,-1,-1,-1,
14'h1944: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,-1,-1,-1,
14'h1945: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,-1,-1,-1,
14'h1946: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,-1,-1,-1,
14'h1947: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,-1,-1,-1,
14'h1950: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,-1,-1,-1,
14'h1951: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,-1,-1,-1,
14'h1952: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,-1,-1,-1,
14'h1953: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,-1,-1,-1,
14'h1954: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,-1,-1,-1,
14'h1955: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,-1,-1,-1,
14'h1956: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,-1,-1,-1,
14'h1957: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //18,19,20,21,22,-1,-1,-1,
14'h1960: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,-1,-1,-1,
14'h1961: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,-1,-1,-1,
14'h1962: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,-1,-1,-1,
14'h1963: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,-1,-1,-1,
14'h1964: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //22,23,24,25,26,-1,-1,-1,
14'h1965: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //22,23,24,25,26,-1,-1,-1,
14'h1966: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //22,23,24,25,26,-1,-1,-1,
14'h1967: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //22,23,24,25,26,-1,-1,-1,
14'h1970: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,-1,-1,-1,
14'h1971: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,-1,-1,-1,
14'h1972: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,-1,-1,-1,
14'h1973: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,-1,-1,-1,
14'h1974: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,-1,-1,-1,
14'h1975: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,-1,-1,-1,
14'h1976: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,-1,-1,-1,
14'h1977: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,-1,-1,-1,
14'h1a00: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,0,1,2,3,
14'h1a01: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 1;   end //0,1,2,3,4,5,6,7,
14'h1a02: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 1; adrVal[7]= 7;   end //0,1,2,3,8,9,10,11,
14'h1a03: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 1; adrVal[4]= 1; adrVal[5]= 1; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,12,13,14,15,
14'h1a04: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,-1,-1,-1,-1,
14'h1a05: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,-1,-1,-1,-1,
14'h1a06: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,-1,-1,-1,-1,
14'h1a07: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,-1,-1,-1,-1,
14'h1a10: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,-1,-1,-1,-1,
14'h1a11: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,-1,-1,-1,-1,
14'h1a12: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,-1,-1,-1,-1,
14'h1a13: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,-1,-1,-1,-1,
14'h1a14: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,-1,-1,-1,-1,
14'h1a15: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,-1,-1,-1,-1,
14'h1a16: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,-1,-1,-1,-1,
14'h1a17: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,-1,-1,-1,-1,
14'h1a20: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h1a21: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h1a22: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h1a23: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h1a24: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h1a25: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h1a26: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h1a27: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,-1,-1,-1,-1,
14'h1a30: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h1a31: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h1a32: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h1a33: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h1a34: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h1a35: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h1a36: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h1a37: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,-1,-1,-1,-1,
14'h1a40: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h1a41: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h1a42: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h1a43: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h1a44: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h1a45: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h1a46: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h1a47: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,-1,-1,-1,-1,
14'h1a50: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h1a51: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h1a52: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h1a53: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h1a54: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h1a55: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h1a56: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h1a57: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,-1,-1,-1,-1,
14'h1a60: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,-1,-1,-1,-1,
14'h1a61: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,-1,-1,-1,-1,
14'h1a62: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,-1,-1,-1,-1,
14'h1a63: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,-1,-1,-1,-1,
14'h1a64: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,-1,-1,-1,-1,
14'h1a65: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,-1,-1,-1,-1,
14'h1a66: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,-1,-1,-1,-1,
14'h1a67: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,-1,-1,-1,-1,
14'h1a70: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,-1,-1,-1,-1,
14'h1a71: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,-1,-1,-1,-1,
14'h1a72: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,-1,-1,-1,-1,
14'h1a73: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,-1,-1,-1,-1,
14'h1a74: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,-1,-1,-1,-1,
14'h1a75: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,-1,-1,-1,-1,
14'h1a76: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,-1,-1,-1,-1,
14'h1a77: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,-1,-1,-1,-1,
14'h1b00: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,-1,-1,
14'h1b01: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,-1,-1,
14'h1b02: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,-1,-1,
14'h1b03: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,-1,-1,
14'h1b04: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,-1,-1,
14'h1b05: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,-1,-1,
14'h1b06: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,-1,-1,
14'h1b07: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,-1,-1,
14'h1b10: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,-1,-1,
14'h1b11: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,-1,-1,
14'h1b12: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,-1,-1,
14'h1b13: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,-1,-1,
14'h1b14: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h1b15: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h1b16: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h1b17: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h1b20: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h1b21: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h1b22: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h1b23: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h1b24: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h1b25: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h1b26: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h1b27: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h1b30: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h1b31: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h1b32: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h1b33: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h1b34: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h1b35: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h1b36: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h1b37: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h1b40: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h1b41: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h1b42: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h1b43: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h1b44: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h1b45: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h1b46: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h1b47: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h1b50: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h1b51: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h1b52: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h1b53: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h1b54: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h1b55: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h1b56: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h1b57: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h1b60: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,-1,-1,
14'h1b61: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,-1,-1,
14'h1b62: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,-1,-1,
14'h1b63: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,-1,-1,
14'h1b64: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,-1,-1,
14'h1b65: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,-1,-1,
14'h1b66: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,-1,-1,
14'h1b67: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,-1,-1,
14'h1b70: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,-1,-1,
14'h1b71: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,-1,-1,
14'h1b72: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,-1,-1,
14'h1b73: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,-1,-1,
14'h1b74: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,-1,-1,
14'h1b75: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,-1,-1,
14'h1b76: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,-1,-1,
14'h1b77: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,-1,-1,
14'h1c00: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,-1,-1,
14'h1c01: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,-1,-1,
14'h1c02: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,-1,-1,
14'h1c03: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,7,-1,-1,
14'h1c04: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,7,-1,-1,
14'h1c05: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,-1,-1,
14'h1c06: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,-1,-1,
14'h1c07: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,-1,-1,
14'h1c10: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,-1,-1,
14'h1c11: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,-1,-1,
14'h1c12: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h1c13: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,11,-1,-1,
14'h1c14: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,11,-1,-1,
14'h1c15: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h1c16: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h1c17: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h1c20: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h1c21: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h1c22: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h1c23: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,-1,-1,
14'h1c24: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,-1,-1,
14'h1c25: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h1c26: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h1c27: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h1c30: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h1c31: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h1c32: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h1c33: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,-1,-1,
14'h1c34: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,-1,-1,
14'h1c35: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h1c36: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h1c37: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h1c40: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h1c41: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h1c42: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h1c43: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,-1,-1,
14'h1c44: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,-1,-1,
14'h1c45: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h1c46: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h1c47: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h1c50: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h1c51: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h1c52: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h1c53: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //22,23,24,25,26,27,-1,-1,
14'h1c54: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //22,23,24,25,26,27,-1,-1,
14'h1c55: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,-1,-1,
14'h1c56: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,-1,-1,
14'h1c57: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,-1,-1,
14'h1c60: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,-1,-1,
14'h1c61: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,-1,-1,
14'h1c62: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,-1,-1,
14'h1c63: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,31,-1,-1,
14'h1c64: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,31,-1,-1,
14'h1c65: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,32,-1,-1,
14'h1c66: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,32,-1,-1,
14'h1c67: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,-1,-1,
14'h1c70: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,-1,-1,
14'h1c71: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,-1,-1,
14'h1c72: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,-1,-1,
14'h1c73: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //30,31,32,33,34,35,-1,-1,
14'h1c74: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //30,31,32,33,34,35,-1,-1,
14'h1c75: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //31,32,33,34,35,36,-1,-1,
14'h1c76: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //31,32,33,34,35,36,-1,-1,
14'h1c77: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //32,33,34,35,36,37,-1,-1,
14'h1d00: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,-1,-1,
14'h1d01: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,-1,-1,
14'h1d02: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,7,-1,-1,
14'h1d03: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,-1,-1,
14'h1d04: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,-1,-1,
14'h1d05: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h1d06: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h1d07: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h1d10: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,-1,-1,
14'h1d11: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,-1,-1,
14'h1d12: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,11,-1,-1,
14'h1d13: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,-1,-1,
14'h1d14: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h1d15: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h1d16: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h1d17: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h1d20: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,-1,-1,
14'h1d21: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,-1,-1,
14'h1d22: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,-1,-1,
14'h1d23: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,-1,-1,
14'h1d24: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h1d25: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h1d26: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h1d27: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h1d30: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,-1,-1,
14'h1d31: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,-1,-1,
14'h1d32: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,-1,-1,
14'h1d33: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,-1,-1,
14'h1d34: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h1d35: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h1d36: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h1d37: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h1d40: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,-1,-1,
14'h1d41: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //17,18,19,20,21,22,-1,-1,
14'h1d42: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,-1,-1,
14'h1d43: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,-1,-1,
14'h1d44: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h1d45: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h1d46: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,-1,-1,
14'h1d47: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,-1,-1,
14'h1d50: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,-1,-1,
14'h1d51: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //21,22,23,24,25,26,-1,-1,
14'h1d52: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //22,23,24,25,26,27,-1,-1,
14'h1d53: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,-1,-1,
14'h1d54: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,-1,-1,
14'h1d55: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,-1,-1,
14'h1d56: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,32,-1,-1,
14'h1d57: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,-1,-1,
14'h1d60: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,-1,-1,
14'h1d61: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,-1,-1,
14'h1d62: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,31,-1,-1,
14'h1d63: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,32,-1,-1,
14'h1d64: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,-1,-1,
14'h1d65: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,-1,-1,
14'h1d66: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //31,32,33,34,35,36,-1,-1,
14'h1d67: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //32,33,34,35,36,37,-1,-1,
14'h1d70: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,-1,-1,
14'h1d71: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,-1,-1,
14'h1d72: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //30,31,32,33,34,35,-1,-1,
14'h1d73: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //31,32,33,34,35,36,-1,-1,
14'h1d74: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //32,33,34,35,36,37,-1,-1,
14'h1d75: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //33,34,35,36,37,38,-1,-1,
14'h1d76: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //35,36,37,38,39,40,-1,-1,
14'h1d77: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //36,37,38,39,40,41,-1,-1,
14'h1e00: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,-1,
14'h1e01: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,7,8,-1,
14'h1e02: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,9,-1,
14'h1e03: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h1e04: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,11,12,-1,
14'h1e05: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h1e06: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h1e07: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h1e10: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,-1,
14'h1e11: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,11,12,-1,
14'h1e12: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h1e13: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h1e14: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h1e15: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h1e16: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h1e17: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h1e20: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h1e21: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h1e22: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h1e23: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h1e24: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h1e25: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h1e26: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,24,-1,
14'h1e27: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h1e30: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h1e31: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h1e32: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h1e33: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h1e34: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,24,-1,
14'h1e35: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h1e36: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //22,23,24,25,26,27,28,-1,
14'h1e37: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,29,-1,
14'h1e40: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h1e41: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,24,-1,
14'h1e42: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h1e43: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,-1,
14'h1e44: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //22,23,24,25,26,27,28,-1,
14'h1e45: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,30,-1,
14'h1e46: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,31,32,-1,
14'h1e47: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,32,33,-1,
14'h1e50: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h1e51: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //22,23,24,25,26,27,28,-1,
14'h1e52: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,29,-1,
14'h1e53: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,31,-1,
14'h1e54: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,31,32,-1,
14'h1e55: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,34,-1,
14'h1e56: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //30,31,32,33,34,35,36,-1,
14'h1e57: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //31,32,33,34,35,36,37,-1,
14'h1e60: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,30,-1,
14'h1e61: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,31,32,-1,
14'h1e62: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,32,33,-1,
14'h1e63: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,35,-1,
14'h1e64: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //30,31,32,33,34,35,36,-1,
14'h1e65: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //32,33,34,35,36,37,38,-1,
14'h1e66: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //34,35,36,37,38,39,40,-1,
14'h1e67: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //35,36,37,38,39,40,41,-1,
14'h1e70: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,34,-1,
14'h1e71: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //30,31,32,33,34,35,36,-1,
14'h1e72: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //31,32,33,34,35,36,37,-1,
14'h1e73: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //33,34,35,36,37,38,39,-1,
14'h1e74: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //34,35,36,37,38,39,40,-1,
14'h1e75: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //36,37,38,39,40,41,42,-1,
14'h1e76: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //38,39,40,41,42,43,44,-1,
14'h1e77: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //39,40,41,42,43,44,45,-1,
14'h1f00: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,-1,
14'h1f01: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //2,3,4,5,6,7,8,-1,
14'h1f02: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,-1,
14'h1f03: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,11,12,-1,
14'h1f04: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h1f05: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h1f06: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h1f07: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h1f10: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,-1,
14'h1f11: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //6,7,8,9,10,11,12,-1,
14'h1f12: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h1f13: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h1f14: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h1f15: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h1f16: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h1f17: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h1f20: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h1f21: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,-1,
14'h1f22: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h1f23: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h1f24: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h1f25: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h1f26: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,-1,
14'h1f27: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,29,-1,
14'h1f30: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h1f31: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,-1,
14'h1f32: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h1f33: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,24,-1,
14'h1f34: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,-1,
14'h1f35: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,29,-1,
14'h1f36: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,31,-1,
14'h1f37: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,32,33,-1,
14'h1f40: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h1f41: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,24,-1,
14'h1f42: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h1f43: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //22,23,24,25,26,27,28,-1,
14'h1f44: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,31,-1,
14'h1f45: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,32,33,-1,
14'h1f46: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,35,-1,
14'h1f47: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //31,32,33,34,35,36,37,-1,
14'h1f50: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h1f51: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //22,23,24,25,26,27,28,-1,
14'h1f52: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,30,-1,
14'h1f53: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,31,32,-1,
14'h1f54: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,35,-1,
14'h1f55: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //31,32,33,34,35,36,37,-1,
14'h1f56: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //33,34,35,36,37,38,39,-1,
14'h1f57: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //35,36,37,38,39,40,41,-1,
14'h1f60: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,30,-1,
14'h1f61: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,31,32,-1,
14'h1f62: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,34,-1,
14'h1f63: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //30,31,32,33,34,35,36,-1,
14'h1f64: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //33,34,35,36,37,38,39,-1,
14'h1f65: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //35,36,37,38,39,40,41,-1,
14'h1f66: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //37,38,39,40,41,42,43,-1,
14'h1f67: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //39,40,41,42,43,44,45,-1,
14'h1f70: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,34,-1,
14'h1f71: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //30,31,32,33,34,35,36,-1,
14'h1f72: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //32,33,34,35,36,37,38,-1,
14'h1f73: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //34,35,36,37,38,39,40,-1,
14'h1f74: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //37,38,39,40,41,42,43,-1,
14'h1f75: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //39,40,41,42,43,44,45,-1,
14'h1f76: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,-1,
14'h1f77: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //43,44,45,46,47,48,49,-1,
14'h2000: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,-1,
14'h2001: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //3,4,5,6,7,8,9,-1,
14'h2002: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,11,-1,
14'h2003: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h2004: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h2005: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h2006: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h2007: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h2010: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,-1,
14'h2011: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,13,-1,
14'h2012: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,-1,
14'h2013: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h2014: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h2015: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h2016: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h2017: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,29,-1,
14'h2020: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,-1,
14'h2021: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,-1,
14'h2022: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,-1,
14'h2023: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h2024: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h2025: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,-1,
14'h2026: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,30,-1,
14'h2027: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,32,33,-1,
14'h2030: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,-1,
14'h2031: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,-1,
14'h2032: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,-1,
14'h2033: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h2034: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,29,-1,
14'h2035: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,31,-1,
14'h2036: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,34,-1,
14'h2037: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //31,32,33,34,35,36,37,-1,
14'h2040: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //16,17,18,19,20,21,22,-1,
14'h2041: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,25,-1,
14'h2042: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,-1,
14'h2043: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,30,-1,
14'h2044: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,32,33,-1,
14'h2045: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,35,-1,
14'h2046: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //32,33,34,35,36,37,38,-1,
14'h2047: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //35,36,37,38,39,40,41,-1,
14'h2050: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //20,21,22,23,24,25,26,-1,
14'h2051: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,29,-1,
14'h2052: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,31,-1,
14'h2053: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,34,-1,
14'h2054: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //31,32,33,34,35,36,37,-1,
14'h2055: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //33,34,35,36,37,38,39,-1,
14'h2056: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //36,37,38,39,40,41,42,-1,
14'h2057: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //39,40,41,42,43,44,45,-1,
14'h2060: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,30,-1,
14'h2061: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,32,33,-1,
14'h2062: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,35,-1,
14'h2063: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //32,33,34,35,36,37,38,-1,
14'h2064: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //35,36,37,38,39,40,41,-1,
14'h2065: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //37,38,39,40,41,42,43,-1,
14'h2066: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //40,41,42,43,44,45,46,-1,
14'h2067: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //43,44,45,46,47,48,49,-1,
14'h2070: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,34,-1,
14'h2071: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //31,32,33,34,35,36,37,-1,
14'h2072: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //33,34,35,36,37,38,39,-1,
14'h2073: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //36,37,38,39,40,41,42,-1,
14'h2074: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //39,40,41,42,43,44,45,-1,
14'h2075: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,-1,
14'h2076: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //44,45,46,47,48,49,50,-1,
14'h2077: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 2; adrVal[6]= 7; adrVal[7]= 7;   end //47,48,49,50,51,52,53,-1,
14'h2100: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //0,1,2,3,4,5,6,7,
14'h2101: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,11,
14'h2102: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //7,8,9,10,11,12,13,14,
14'h2103: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //10,11,12,13,14,15,16,17,
14'h2104: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,20,
14'h2105: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,24,
14'h2106: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //20,21,22,23,24,25,26,27,
14'h2107: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,29,30,
14'h2110: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //4,5,6,7,8,9,10,11,
14'h2111: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,15,
14'h2112: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //11,12,13,14,15,16,17,18,
14'h2113: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //14,15,16,17,18,19,20,21,
14'h2114: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,24,
14'h2115: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,28,
14'h2116: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,30,31,
14'h2117: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,32,33,34,
14'h2120: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //8,9,10,11,12,13,14,15,
14'h2121: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,19,
14'h2122: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //15,16,17,18,19,20,21,22,
14'h2123: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //18,19,20,21,22,23,24,25,
14'h2124: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,28,
14'h2125: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,31,32,
14'h2126: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,34,35,
14'h2127: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //31,32,33,34,35,36,37,38,
14'h2130: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //12,13,14,15,16,17,18,19,
14'h2131: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //16,17,18,19,20,21,22,23,
14'h2132: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //19,20,21,22,23,24,25,26,
14'h2133: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //22,23,24,25,26,27,28,29,
14'h2134: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,31,32,
14'h2135: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,35,36,
14'h2136: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //32,33,34,35,36,37,38,39,
14'h2137: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //35,36,37,38,39,40,41,42,
14'h2140: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //16,17,18,19,20,21,22,23,
14'h2141: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //20,21,22,23,24,25,26,27,
14'h2142: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //23,24,25,26,27,28,29,30,
14'h2143: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //26,27,28,29,30,31,32,33,
14'h2144: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,35,36,
14'h2145: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //33,34,35,36,37,38,39,40,
14'h2146: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //36,37,38,39,40,41,42,43,
14'h2147: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //39,40,41,42,43,44,45,46,
14'h2150: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //20,21,22,23,24,25,26,27,
14'h2151: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,30,31,
14'h2152: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //27,28,29,30,31,32,33,34,
14'h2153: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //30,31,32,33,34,35,36,37,
14'h2154: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //33,34,35,36,37,38,39,40,
14'h2155: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //37,38,39,40,41,42,43,44,
14'h2156: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //40,41,42,43,44,45,46,47,
14'h2157: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //43,44,45,46,47,48,49,50,
14'h2160: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //24,25,26,27,28,29,30,31,
14'h2161: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,34,35,
14'h2162: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //31,32,33,34,35,36,37,38,
14'h2163: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //34,35,36,37,38,39,40,41,
14'h2164: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //37,38,39,40,41,42,43,44,
14'h2165: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,48,
14'h2166: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 2; adrVal[6]= 7; adrVal[7]= 7;   end //44,45,46,47,48,49,50,51,
14'h2167: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 2; adrVal[6]= 7; adrVal[7]= 7;   end //47,48,49,50,51,52,53,54,
14'h2170: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //28,29,30,31,32,33,34,35,
14'h2171: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //32,33,34,35,36,37,38,39,
14'h2172: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //35,36,37,38,39,40,41,42,
14'h2173: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //38,39,40,41,42,43,44,45,
14'h2174: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,48,
14'h2175: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 2; adrVal[6]= 7; adrVal[7]= 7;   end //45,46,47,48,49,50,51,52,
14'h2176: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 2; adrVal[6]= 2; adrVal[7]= 7;   end //48,49,50,51,52,53,54,55,
14'h2177: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 2; adrVal[5]= 2; adrVal[6]= 2; adrVal[7]= 7;   end //51,52,53,54,55,56,57,58,
14'h2200: begin  adrVal[0]= 0; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //1,2,3,4,5,6,7,8,
14'h2201: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,11,12,
14'h2202: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,16,
14'h2203: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,20,
14'h2204: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,24,
14'h2205: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,28,
14'h2206: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,31,32,
14'h2207: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,35,36,
14'h2210: begin  adrVal[0]= 7; adrVal[1]= 0; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //5,6,7,8,9,10,11,12,
14'h2211: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,16,
14'h2212: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,20,
14'h2213: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,24,
14'h2214: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,28,
14'h2215: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,31,32,
14'h2216: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,35,36,
14'h2217: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //33,34,35,36,37,38,39,40,
14'h2220: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 0; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //9,10,11,12,13,14,15,16,
14'h2221: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,20,
14'h2222: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,24,
14'h2223: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,28,
14'h2224: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,31,32,
14'h2225: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,35,36,
14'h2226: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //33,34,35,36,37,38,39,40,
14'h2227: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //37,38,39,40,41,42,43,44,
14'h2230: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 0; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 7; adrVal[7]= 7;   end //13,14,15,16,17,18,19,20,
14'h2231: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,24,
14'h2232: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,28,
14'h2233: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,31,32,
14'h2234: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,35,36,
14'h2235: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //33,34,35,36,37,38,39,40,
14'h2236: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //37,38,39,40,41,42,43,44,
14'h2237: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,48,
14'h2240: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 0; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 7;   end //17,18,19,20,21,22,23,24,
14'h2241: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,28,
14'h2242: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,31,32,
14'h2243: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,35,36,
14'h2244: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //33,34,35,36,37,38,39,40,
14'h2245: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //37,38,39,40,41,42,43,44,
14'h2246: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,48,
14'h2247: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 2; adrVal[6]= 7; adrVal[7]= 7;   end //45,46,47,48,49,50,51,52,
14'h2250: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 0; adrVal[6]= 0; adrVal[7]= 0;   end //21,22,23,24,25,26,27,28,
14'h2251: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,31,32,
14'h2252: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,35,36,
14'h2253: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //33,34,35,36,37,38,39,40,
14'h2254: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //37,38,39,40,41,42,43,44,
14'h2255: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,48,
14'h2256: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 2; adrVal[6]= 7; adrVal[7]= 7;   end //45,46,47,48,49,50,51,52,
14'h2257: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 2; adrVal[5]= 2; adrVal[6]= 2; adrVal[7]= 7;   end //49,50,51,52,53,54,55,56,
14'h2260: begin  adrVal[0]= 2; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 0; adrVal[7]= 0;   end //25,26,27,28,29,30,31,32,
14'h2261: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,35,36,
14'h2262: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //33,34,35,36,37,38,39,40,
14'h2263: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //37,38,39,40,41,42,43,44,
14'h2264: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,48,
14'h2265: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 2; adrVal[6]= 7; adrVal[7]= 7;   end //45,46,47,48,49,50,51,52,
14'h2266: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 2; adrVal[5]= 2; adrVal[6]= 2; adrVal[7]= 7;   end //49,50,51,52,53,54,55,56,
14'h2267: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 2; adrVal[6]= 2; adrVal[7]= 2;   end //53,54,55,56,57,58,59,60,
14'h2270: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 0;   end //29,30,31,32,33,34,35,36,
14'h2271: begin  adrVal[0]= 2; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //33,34,35,36,37,38,39,40,
14'h2272: begin  adrVal[0]= 7; adrVal[1]= 2; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //37,38,39,40,41,42,43,44,
14'h2273: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 2; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end //41,42,43,44,45,46,47,48,
14'h2274: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 2; adrVal[4]= 2; adrVal[5]= 2; adrVal[6]= 7; adrVal[7]= 7;   end //45,46,47,48,49,50,51,52,
14'h2275: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 2; adrVal[5]= 2; adrVal[6]= 2; adrVal[7]= 7;   end //49,50,51,52,53,54,55,56,
14'h2276: begin  adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 2; adrVal[6]= 2; adrVal[7]= 2;   end //53,54,55,56,57,58,59,60,
14'h2277: begin  adrVal[0]= 4; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 2; adrVal[7]= 2;   end //57,58,59,60,61,62,63,64,



default: begin adrVal[0]= 7; adrVal[1]= 7; adrVal[2]= 7; adrVal[3]= 7; adrVal[4]= 7; adrVal[5]= 7; adrVal[6]= 7; adrVal[7]= 7;   end 

endcase
end	// end of if(preStage[2] == 1'b1)
endcase
end
endmodule
