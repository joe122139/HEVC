`timescale 1ns/1ps
module intra_refPosGen(
	mode,			//i
	X,				//i
	Y,
	ref_pos,   //o
	ref_TLADflag  //o
	,preStage
	,tuSize
);


input [5:0] mode;
input [2:0] X;
input [2:0] Y;
input [3:0] preStage; 
input [2:0] tuSize;
  

output reg [47:0] ref_pos;
output reg [15:0] ref_TLADflag;	//0 top,  1 left, 2 top_left , 

  
reg [5:0] refPos[7:0];		//dp
reg [1:0] refFlag[7:0];
 

generate
  genvar i;
    for(i=0;i<8;i=i+1)  begin:xi
    always @(*) begin
    //  ref_pos[(55-7*i):(49-7*i)] = refPos[i];
      ref_pos[(47-6*i):(42-6*i)] = refPos[i];
	  ref_TLADflag[(15-2*i):(14-2*i)] = refFlag[i];
    end
  end
endgenerate


always@ (*) begin
	refPos[0]=0; refFlag[0]=0; refPos[1]=0; refFlag[1]=0; refPos[2]=0; refFlag[2]=0; refPos[3]=0; refFlag[3]=0; refPos[4]=0; refFlag[4]=0; refPos[5]=0; refFlag[5]=0; refPos[6]=0; refFlag[6]=0; refPos[7]=0; refFlag[7]=0; 
	if (preStage== 0 && tuSize== 4)  begin 
		refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=18; refFlag[7]=0; 
	end
	

	else if (preStage== 2)  begin 
		refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=34; refFlag[6]=1; refPos[7]=34; refFlag[7]=1; 
	end

	else if(preStage == 3) begin 
		refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=34; refFlag[6]=0; refPos[7]=34; refFlag[7]=0; 

	end 
	else 

 case({mode,1'b0,X,1'b0,Y})

14'h 000: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h 001: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 002: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 003: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 004: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 005: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 006: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 007: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 010:
	if(tuSize==3'd3)
		begin refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;end
	else
		begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 011: 
		if(tuSize==3'd3)
			begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
		else begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 012: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 013: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 014: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 015: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 016: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 017: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 020: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 021: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 022: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 023: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 024: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 025: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 026: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 027: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 030: 
	if(tuSize==3'd4) 
		begin refPos[0]=1; refFlag[0]=-1; refPos[1]=1; refFlag[1]=-1; refPos[2]=1; refFlag[2]=-1; refPos[3]=1; refFlag[3]=-1; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
	else 
		begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 031: if(tuSize==3'd4)  
		begin refPos[0]=1; refFlag[0]=-1; refPos[1]=1; refFlag[1]=-1; refPos[2]=1; refFlag[2]=-1; refPos[3]=1; refFlag[3]=-1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
	else 
		begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
		
14'h 032: 
	if(tuSize==3'd4) 
		begin refPos[0]=1; refFlag[0]=-1; refPos[1]=1; refFlag[1]=-1; refPos[2]=1; refFlag[2]=-1; refPos[3]=1; refFlag[3]=-1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
	else
		begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 033: 
	if(tuSize==3'd4) 
		begin refPos[0]=15; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
	else
		begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 034: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 035: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 036: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 037: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 040: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 041: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 042: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 043: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 044: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 045: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 046: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 047: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 050: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 051: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 052: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 053: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 054: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 055: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 056: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 057: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 060: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 061: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 062: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 063: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 064: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 065: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 066: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 067: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 070: if(tuSize== 5) 
	begin refPos[0]=1; refFlag[0]=-1; refPos[1]=1; refFlag[1]=-1; refPos[2]=1; refFlag[2]=-1; refPos[3]=1; refFlag[3]=-1; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
	else
	begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 

14'h 071: if(tuSize== 5) 
		begin refPos[0]=1; refFlag[0]=-1; refPos[1]=1; refFlag[1]=-1; refPos[2]=1; refFlag[2]=-1; refPos[3]=1; refFlag[3]=-1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
	else begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 072: if(tuSize== 5) 
			begin refPos[0]=1; refFlag[0]=-1; refPos[1]=1; refFlag[1]=-1; refPos[2]=1; refFlag[2]=-1; refPos[3]=1; refFlag[3]=-1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
		else
			begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 073: if(tuSize== 5) 
			begin refPos[0]=1; refFlag[0]=-1; refPos[1]=1; refFlag[1]=-1; refPos[2]=1; refFlag[2]=-1; refPos[3]=1; refFlag[3]=-1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
		else begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 074: if(tuSize== 5)
			begin refPos[0]=1; refFlag[0]=-1; refPos[1]=1; refFlag[1]=-1; refPos[2]=1; refFlag[2]=-1; refPos[3]=1; refFlag[3]=-1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=19; refFlag[7]=1;  end 
		else
			begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 075: if(tuSize== 5)
			begin refPos[0]=1; refFlag[0]=-1; refPos[1]=1; refFlag[1]=-1; refPos[2]=1; refFlag[2]=-1; refPos[3]=1; refFlag[3]=-1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=23; refFlag[7]=1;  end 
		else
			begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 076: if(tuSize== 5)
			begin refPos[0]=1; refFlag[0]=-1; refPos[1]=1; refFlag[1]=-1; refPos[2]=1; refFlag[2]=-1; refPos[3]=1; refFlag[3]=-1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=27; refFlag[7]=1;  end 
		else 
			begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 077: if(tuSize== 5) 
			begin refPos[0]=1; refFlag[0]=-1; refPos[1]=1; refFlag[1]=-1; refPos[2]=1; refFlag[2]=-1; refPos[3]=1; refFlag[3]=-1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=31; refFlag[7]=1;  end 
		else begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h 100: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h 101: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h 102: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h 103: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
14'h 104: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=19; refFlag[7]=1;  end 
14'h 105: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=23; refFlag[7]=1;  end 
14'h 106: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=27; refFlag[7]=1;  end 
14'h 107: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=31; refFlag[7]=1;  end 
14'h 110: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h 111: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h 112: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h 113: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
14'h 114: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=19; refFlag[7]=1;  end 
14'h 115: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=23; refFlag[7]=1;  end 
14'h 116: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=27; refFlag[7]=1;  end 
14'h 117: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=31; refFlag[7]=1;  end 
14'h 120: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h 121: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h 122: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h 123: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
14'h 124: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=19; refFlag[7]=1;  end 
14'h 125: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=23; refFlag[7]=1;  end 
14'h 126: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=27; refFlag[7]=1;  end 
14'h 127: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=31; refFlag[7]=1;  end 
14'h 130: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h 131: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h 132: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h 133: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
14'h 134: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=19; refFlag[7]=1;  end 
14'h 135: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=23; refFlag[7]=1;  end 
14'h 136: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=27; refFlag[7]=1;  end 
14'h 137: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=31; refFlag[7]=1;  end 
14'h 140: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h 141: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h 142: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h 143: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
14'h 144: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=19; refFlag[7]=1;  end 
14'h 145: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=23; refFlag[7]=1;  end 
14'h 146: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=27; refFlag[7]=1;  end 
14'h 147: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=31; refFlag[7]=1;  end 
14'h 150: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h 151: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h 152: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h 153: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
14'h 154: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=19; refFlag[7]=1;  end 
14'h 155: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=23; refFlag[7]=1;  end 
14'h 156: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=27; refFlag[7]=1;  end 
14'h 157: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=31; refFlag[7]=1;  end 
14'h 160: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h 161: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h 162: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h 163: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
14'h 164: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=19; refFlag[7]=1;  end 
14'h 165: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=23; refFlag[7]=1;  end 
14'h 166: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=27; refFlag[7]=1;  end 
14'h 167: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=31; refFlag[7]=1;  end 
14'h 170: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h 171: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h 172: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h 173: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
14'h 174: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=19; refFlag[7]=1;  end 
14'h 175: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=23; refFlag[7]=1;  end 
14'h 176: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=27; refFlag[7]=1;  end 
14'h 177: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=31; refFlag[7]=1;  end 
14'h 200: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=7; refFlag[6]=1; if(tuSize!=2) refPos[7]=8; else refPos[7]=7; refFlag[7]=1;  end 
14'h 201: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=12; refFlag[7]=1;  end 
14'h 202: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=15; refFlag[6]=1; refPos[7]=16; refFlag[7]=1;  end 
14'h 203: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=20; refFlag[7]=1;  end 
14'h 204: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=24; refFlag[7]=1;  end 
14'h 205: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=28; refFlag[7]=1;  end 
14'h 206: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=31; refFlag[6]=1; refPos[7]=32; refFlag[7]=1;  end 
14'h 207: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=35; refFlag[6]=1; refPos[7]=36; refFlag[7]=1;  end 
14'h 210: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=12; refFlag[7]=1;  end 
14'h 211: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=15; refFlag[6]=1; if(tuSize!=3)refPos[7]=16; else refPos[7]=15;  refFlag[7]=1;  end 
14'h 212: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=20; refFlag[7]=1;  end 
14'h 213: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=24; refFlag[7]=1;  end 
14'h 214: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=28; refFlag[7]=1;  end 
14'h 215: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=31; refFlag[6]=1; refPos[7]=32; refFlag[7]=1;  end 
14'h 216: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=35; refFlag[6]=1; refPos[7]=36; refFlag[7]=1;  end 
14'h 217: begin refPos[0]=33; refFlag[0]=1; refPos[1]=34; refFlag[1]=1; refPos[2]=35; refFlag[2]=1; refPos[3]=36; refFlag[3]=1; refPos[4]=37; refFlag[4]=1; refPos[5]=38; refFlag[5]=1; refPos[6]=39; refFlag[6]=1; refPos[7]=40; refFlag[7]=1;  end 
14'h 220: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=15; refFlag[6]=1; refPos[7]=16; refFlag[7]=1;  end 
14'h 221: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=20; refFlag[7]=1;  end 
14'h 222: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=24; refFlag[7]=1;  end 
14'h 223: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=28; refFlag[7]=1;  end 
14'h 224: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=31; refFlag[6]=1; refPos[7]=32; refFlag[7]=1;  end 
14'h 225: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=35; refFlag[6]=1; refPos[7]=36; refFlag[7]=1;  end 
14'h 226: begin refPos[0]=33; refFlag[0]=1; refPos[1]=34; refFlag[1]=1; refPos[2]=35; refFlag[2]=1; refPos[3]=36; refFlag[3]=1; refPos[4]=37; refFlag[4]=1; refPos[5]=38; refFlag[5]=1; refPos[6]=39; refFlag[6]=1; refPos[7]=40; refFlag[7]=1;  end 
14'h 227: begin refPos[0]=37; refFlag[0]=1; refPos[1]=38; refFlag[1]=1; refPos[2]=39; refFlag[2]=1; refPos[3]=40; refFlag[3]=1; refPos[4]=41; refFlag[4]=1; refPos[5]=42; refFlag[5]=1; refPos[6]=43; refFlag[6]=1; refPos[7]=44; refFlag[7]=1;  end 
14'h 230: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=20; refFlag[7]=1;  end 
14'h 231: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=24; refFlag[7]=1;  end 
14'h 232: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=28; refFlag[7]=1;  end 
14'h 233: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=31; refFlag[6]=1; if(tuSize!=4) refPos[7]=32; else refPos[7]=31; refFlag[7]=1;  end 
14'h 234: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=35; refFlag[6]=1; refPos[7]=36; refFlag[7]=1;  end 
14'h 235: begin refPos[0]=33; refFlag[0]=1; refPos[1]=34; refFlag[1]=1; refPos[2]=35; refFlag[2]=1; refPos[3]=36; refFlag[3]=1; refPos[4]=37; refFlag[4]=1; refPos[5]=38; refFlag[5]=1; refPos[6]=39; refFlag[6]=1; refPos[7]=40; refFlag[7]=1;  end 
14'h 236: begin refPos[0]=37; refFlag[0]=1; refPos[1]=38; refFlag[1]=1; refPos[2]=39; refFlag[2]=1; refPos[3]=40; refFlag[3]=1; refPos[4]=41; refFlag[4]=1; refPos[5]=42; refFlag[5]=1; refPos[6]=43; refFlag[6]=1; refPos[7]=44; refFlag[7]=1;  end 
14'h 237: begin refPos[0]=41; refFlag[0]=1; refPos[1]=42; refFlag[1]=1; refPos[2]=43; refFlag[2]=1; refPos[3]=44; refFlag[3]=1; refPos[4]=45; refFlag[4]=1; refPos[5]=46; refFlag[5]=1; refPos[6]=47; refFlag[6]=1; refPos[7]=48; refFlag[7]=1;  end 
14'h 240: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=24; refFlag[7]=1;  end 
14'h 241: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=28; refFlag[7]=1;  end 
14'h 242: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=31; refFlag[6]=1; refPos[7]=32; refFlag[7]=1;  end 
14'h 243: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=35; refFlag[6]=1; refPos[7]=36; refFlag[7]=1;  end 
14'h 244: begin refPos[0]=33; refFlag[0]=1; refPos[1]=34; refFlag[1]=1; refPos[2]=35; refFlag[2]=1; refPos[3]=36; refFlag[3]=1; refPos[4]=37; refFlag[4]=1; refPos[5]=38; refFlag[5]=1; refPos[6]=39; refFlag[6]=1; refPos[7]=40; refFlag[7]=1;  end 
14'h 245: begin refPos[0]=37; refFlag[0]=1; refPos[1]=38; refFlag[1]=1; refPos[2]=39; refFlag[2]=1; refPos[3]=40; refFlag[3]=1; refPos[4]=41; refFlag[4]=1; refPos[5]=42; refFlag[5]=1; refPos[6]=43; refFlag[6]=1; refPos[7]=44; refFlag[7]=1;  end 
14'h 246: begin refPos[0]=41; refFlag[0]=1; refPos[1]=42; refFlag[1]=1; refPos[2]=43; refFlag[2]=1; refPos[3]=44; refFlag[3]=1; refPos[4]=45; refFlag[4]=1; refPos[5]=46; refFlag[5]=1; refPos[6]=47; refFlag[6]=1; refPos[7]=48; refFlag[7]=1;  end 
14'h 247: begin refPos[0]=45; refFlag[0]=1; refPos[1]=46; refFlag[1]=1; refPos[2]=47; refFlag[2]=1; refPos[3]=48; refFlag[3]=1; refPos[4]=49; refFlag[4]=1; refPos[5]=50; refFlag[5]=1; refPos[6]=51; refFlag[6]=1; refPos[7]=52; refFlag[7]=1;  end 
14'h 250: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=28; refFlag[7]=1;  end 
14'h 251: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=31; refFlag[6]=1; refPos[7]=32; refFlag[7]=1;  end 
14'h 252: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=35; refFlag[6]=1; refPos[7]=36; refFlag[7]=1;  end 
14'h 253: begin refPos[0]=33; refFlag[0]=1; refPos[1]=34; refFlag[1]=1; refPos[2]=35; refFlag[2]=1; refPos[3]=36; refFlag[3]=1; refPos[4]=37; refFlag[4]=1; refPos[5]=38; refFlag[5]=1; refPos[6]=39; refFlag[6]=1; refPos[7]=40; refFlag[7]=1;  end 
14'h 254: begin refPos[0]=37; refFlag[0]=1; refPos[1]=38; refFlag[1]=1; refPos[2]=39; refFlag[2]=1; refPos[3]=40; refFlag[3]=1; refPos[4]=41; refFlag[4]=1; refPos[5]=42; refFlag[5]=1; refPos[6]=43; refFlag[6]=1; refPos[7]=44; refFlag[7]=1;  end 
14'h 255: begin refPos[0]=41; refFlag[0]=1; refPos[1]=42; refFlag[1]=1; refPos[2]=43; refFlag[2]=1; refPos[3]=44; refFlag[3]=1; refPos[4]=45; refFlag[4]=1; refPos[5]=46; refFlag[5]=1; refPos[6]=47; refFlag[6]=1; refPos[7]=48; refFlag[7]=1;  end 
14'h 256: begin refPos[0]=45; refFlag[0]=1; refPos[1]=46; refFlag[1]=1; refPos[2]=47; refFlag[2]=1; refPos[3]=48; refFlag[3]=1; refPos[4]=49; refFlag[4]=1; refPos[5]=50; refFlag[5]=1; refPos[6]=51; refFlag[6]=1; refPos[7]=52; refFlag[7]=1;  end 
14'h 257: begin refPos[0]=49; refFlag[0]=1; refPos[1]=50; refFlag[1]=1; refPos[2]=51; refFlag[2]=1; refPos[3]=52; refFlag[3]=1; refPos[4]=53; refFlag[4]=1; refPos[5]=54; refFlag[5]=1; refPos[6]=55; refFlag[6]=1; refPos[7]=56; refFlag[7]=1;  end 
14'h 260: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=31; refFlag[6]=1; refPos[7]=32; refFlag[7]=1;  end 
14'h 261: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=35; refFlag[6]=1; refPos[7]=36; refFlag[7]=1;  end 
14'h 262: begin refPos[0]=33; refFlag[0]=1; refPos[1]=34; refFlag[1]=1; refPos[2]=35; refFlag[2]=1; refPos[3]=36; refFlag[3]=1; refPos[4]=37; refFlag[4]=1; refPos[5]=38; refFlag[5]=1; refPos[6]=39; refFlag[6]=1; refPos[7]=40; refFlag[7]=1;  end 
14'h 263: begin refPos[0]=37; refFlag[0]=1; refPos[1]=38; refFlag[1]=1; refPos[2]=39; refFlag[2]=1; refPos[3]=40; refFlag[3]=1; refPos[4]=41; refFlag[4]=1; refPos[5]=42; refFlag[5]=1; refPos[6]=43; refFlag[6]=1; refPos[7]=44; refFlag[7]=1;  end 
14'h 264: begin refPos[0]=41; refFlag[0]=1; refPos[1]=42; refFlag[1]=1; refPos[2]=43; refFlag[2]=1; refPos[3]=44; refFlag[3]=1; refPos[4]=45; refFlag[4]=1; refPos[5]=46; refFlag[5]=1; refPos[6]=47; refFlag[6]=1; refPos[7]=48; refFlag[7]=1;  end 
14'h 265: begin refPos[0]=45; refFlag[0]=1; refPos[1]=46; refFlag[1]=1; refPos[2]=47; refFlag[2]=1; refPos[3]=48; refFlag[3]=1; refPos[4]=49; refFlag[4]=1; refPos[5]=50; refFlag[5]=1; refPos[6]=51; refFlag[6]=1; refPos[7]=52; refFlag[7]=1;  end 
14'h 266: begin refPos[0]=49; refFlag[0]=1; refPos[1]=50; refFlag[1]=1; refPos[2]=51; refFlag[2]=1; refPos[3]=52; refFlag[3]=1; refPos[4]=53; refFlag[4]=1; refPos[5]=54; refFlag[5]=1; refPos[6]=55; refFlag[6]=1; refPos[7]=56; refFlag[7]=1;  end 
14'h 267: begin refPos[0]=53; refFlag[0]=1; refPos[1]=54; refFlag[1]=1; refPos[2]=55; refFlag[2]=1; refPos[3]=56; refFlag[3]=1; refPos[4]=57; refFlag[4]=1; refPos[5]=58; refFlag[5]=1; refPos[6]=59; refFlag[6]=1; refPos[7]=60; refFlag[7]=1;  end 
14'h 270: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=35; refFlag[6]=1; refPos[7]=36; refFlag[7]=1;  end 
14'h 271: begin refPos[0]=33; refFlag[0]=1; refPos[1]=34; refFlag[1]=1; refPos[2]=35; refFlag[2]=1; refPos[3]=36; refFlag[3]=1; refPos[4]=37; refFlag[4]=1; refPos[5]=38; refFlag[5]=1; refPos[6]=39; refFlag[6]=1; refPos[7]=40; refFlag[7]=1;  end 
14'h 272: begin refPos[0]=37; refFlag[0]=1; refPos[1]=38; refFlag[1]=1; refPos[2]=39; refFlag[2]=1; refPos[3]=40; refFlag[3]=1; refPos[4]=41; refFlag[4]=1; refPos[5]=42; refFlag[5]=1; refPos[6]=43; refFlag[6]=1; refPos[7]=44; refFlag[7]=1;  end 
14'h 273: begin refPos[0]=41; refFlag[0]=1; refPos[1]=42; refFlag[1]=1; refPos[2]=43; refFlag[2]=1; refPos[3]=44; refFlag[3]=1; refPos[4]=45; refFlag[4]=1; refPos[5]=46; refFlag[5]=1; refPos[6]=47; refFlag[6]=1; refPos[7]=48; refFlag[7]=1;  end 
14'h 274: begin refPos[0]=45; refFlag[0]=1; refPos[1]=46; refFlag[1]=1; refPos[2]=47; refFlag[2]=1; refPos[3]=48; refFlag[3]=1; refPos[4]=49; refFlag[4]=1; refPos[5]=50; refFlag[5]=1; refPos[6]=51; refFlag[6]=1; refPos[7]=52; refFlag[7]=1;  end 
14'h 275: begin refPos[0]=49; refFlag[0]=1; refPos[1]=50; refFlag[1]=1; refPos[2]=51; refFlag[2]=1; refPos[3]=52; refFlag[3]=1; refPos[4]=53; refFlag[4]=1; refPos[5]=54; refFlag[5]=1; refPos[6]=55; refFlag[6]=1; refPos[7]=56; refFlag[7]=1;  end 
14'h 276: begin refPos[0]=53; refFlag[0]=1; refPos[1]=54; refFlag[1]=1; refPos[2]=55; refFlag[2]=1; refPos[3]=56; refFlag[3]=1; refPos[4]=57; refFlag[4]=1; refPos[5]=58; refFlag[5]=1; refPos[6]=59; refFlag[6]=1; refPos[7]=60; refFlag[7]=1;  end 
14'h 277: begin refPos[0]=57; refFlag[0]=1; refPos[1]=58; refFlag[1]=1; refPos[2]=59; refFlag[2]=1; refPos[3]=60; refFlag[3]=1; refPos[4]=61; refFlag[4]=1; refPos[5]=62; refFlag[5]=1; refPos[6]=63; refFlag[6]=1; refPos[7]=63; refFlag[7]=1;  end 
14'h 300: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h 301: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h 302: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=13; refFlag[6]=1; refPos[7]=14; refFlag[7]=1;  end 
14'h 303: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=16; refFlag[6]=1; refPos[7]=17; refFlag[7]=1;  end 
14'h 304: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=20; refFlag[7]=1;  end 
14'h 305: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=24; refFlag[7]=1;  end 
14'h 306: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=27; refFlag[7]=1;  end 
14'h 307: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=29; refFlag[6]=1; refPos[7]=30; refFlag[7]=1;  end 
14'h 310: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h 311: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
14'h 312: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=18; refFlag[7]=1;  end 
14'h 313: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=20; refFlag[6]=1; refPos[7]=21; refFlag[7]=1;  end 
14'h 314: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=24; refFlag[7]=1;  end 
14'h 315: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=28; refFlag[7]=1;  end 
14'h 316: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=31; refFlag[7]=1;  end 
14'h 317: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=32; refFlag[5]=1; refPos[6]=33; refFlag[6]=1; refPos[7]=34; refFlag[7]=1;  end 
14'h 320: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
14'h 321: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=19; refFlag[7]=1;  end 
14'h 322: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=21; refFlag[6]=1; refPos[7]=22; refFlag[7]=1;  end 
14'h 323: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=24; refFlag[6]=1; refPos[7]=25; refFlag[7]=1;  end 
14'h 324: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=28; refFlag[7]=1;  end 
14'h 325: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=31; refFlag[6]=1; refPos[7]=32; refFlag[7]=1;  end 
14'h 326: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=34; refFlag[6]=1; refPos[7]=35; refFlag[7]=1;  end 
14'h 327: begin refPos[0]=31; refFlag[0]=1; refPos[1]=32; refFlag[1]=1; refPos[2]=33; refFlag[2]=1; refPos[3]=34; refFlag[3]=1; refPos[4]=35; refFlag[4]=1; refPos[5]=36; refFlag[5]=1; refPos[6]=37; refFlag[6]=1; refPos[7]=38; refFlag[7]=1;  end 
14'h 330: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=19; refFlag[7]=1;  end 
14'h 331: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=23; refFlag[7]=1;  end 
14'h 332: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=25; refFlag[6]=1; refPos[7]=26; refFlag[7]=1;  end 
14'h 333: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=27; refFlag[5]=1; refPos[6]=28; refFlag[6]=1; refPos[7]=29; refFlag[7]=1;  end 
14'h 334: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=31; refFlag[6]=1; refPos[7]=32; refFlag[7]=1;  end 
14'h 335: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=35; refFlag[6]=1; refPos[7]=36; refFlag[7]=1;  end 
14'h 336: begin refPos[0]=32; refFlag[0]=1; refPos[1]=33; refFlag[1]=1; refPos[2]=34; refFlag[2]=1; refPos[3]=35; refFlag[3]=1; refPos[4]=36; refFlag[4]=1; refPos[5]=37; refFlag[5]=1; refPos[6]=38; refFlag[6]=1; refPos[7]=39; refFlag[7]=1;  end 
14'h 337: begin refPos[0]=35; refFlag[0]=1; refPos[1]=36; refFlag[1]=1; refPos[2]=37; refFlag[2]=1; refPos[3]=38; refFlag[3]=1; refPos[4]=39; refFlag[4]=1; refPos[5]=40; refFlag[5]=1; refPos[6]=41; refFlag[6]=1; refPos[7]=42; refFlag[7]=1;  end 
14'h 340: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=23; refFlag[7]=1;  end 
14'h 341: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=27; refFlag[7]=1;  end 
14'h 342: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=29; refFlag[6]=1; refPos[7]=30; refFlag[7]=1;  end 
14'h 343: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=31; refFlag[5]=1; refPos[6]=32; refFlag[6]=1; refPos[7]=33; refFlag[7]=1;  end 
14'h 344: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=35; refFlag[6]=1; refPos[7]=36; refFlag[7]=1;  end 
14'h 345: begin refPos[0]=33; refFlag[0]=1; refPos[1]=34; refFlag[1]=1; refPos[2]=35; refFlag[2]=1; refPos[3]=36; refFlag[3]=1; refPos[4]=37; refFlag[4]=1; refPos[5]=38; refFlag[5]=1; refPos[6]=39; refFlag[6]=1; refPos[7]=40; refFlag[7]=1;  end 
14'h 346: begin refPos[0]=36; refFlag[0]=1; refPos[1]=37; refFlag[1]=1; refPos[2]=38; refFlag[2]=1; refPos[3]=39; refFlag[3]=1; refPos[4]=40; refFlag[4]=1; refPos[5]=41; refFlag[5]=1; refPos[6]=42; refFlag[6]=1; refPos[7]=43; refFlag[7]=1;  end 
14'h 347: begin refPos[0]=39; refFlag[0]=1; refPos[1]=40; refFlag[1]=1; refPos[2]=41; refFlag[2]=1; refPos[3]=42; refFlag[3]=1; refPos[4]=43; refFlag[4]=1; refPos[5]=44; refFlag[5]=1; refPos[6]=45; refFlag[6]=1; refPos[7]=46; refFlag[7]=1;  end 
14'h 350: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=27; refFlag[7]=1;  end 
14'h 351: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=31; refFlag[7]=1;  end 
14'h 352: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=32; refFlag[5]=1; refPos[6]=33; refFlag[6]=1; refPos[7]=34; refFlag[7]=1;  end 
14'h 353: begin refPos[0]=30; refFlag[0]=1; refPos[1]=31; refFlag[1]=1; refPos[2]=32; refFlag[2]=1; refPos[3]=33; refFlag[3]=1; refPos[4]=34; refFlag[4]=1; refPos[5]=35; refFlag[5]=1; refPos[6]=36; refFlag[6]=1; refPos[7]=37; refFlag[7]=1;  end 
14'h 354: begin refPos[0]=33; refFlag[0]=1; refPos[1]=34; refFlag[1]=1; refPos[2]=35; refFlag[2]=1; refPos[3]=36; refFlag[3]=1; refPos[4]=37; refFlag[4]=1; refPos[5]=38; refFlag[5]=1; refPos[6]=39; refFlag[6]=1; refPos[7]=40; refFlag[7]=1;  end 
14'h 355: begin refPos[0]=37; refFlag[0]=1; refPos[1]=38; refFlag[1]=1; refPos[2]=39; refFlag[2]=1; refPos[3]=40; refFlag[3]=1; refPos[4]=41; refFlag[4]=1; refPos[5]=42; refFlag[5]=1; refPos[6]=43; refFlag[6]=1; refPos[7]=44; refFlag[7]=1;  end 
14'h 356: begin refPos[0]=40; refFlag[0]=1; refPos[1]=41; refFlag[1]=1; refPos[2]=42; refFlag[2]=1; refPos[3]=43; refFlag[3]=1; refPos[4]=44; refFlag[4]=1; refPos[5]=45; refFlag[5]=1; refPos[6]=46; refFlag[6]=1; refPos[7]=47; refFlag[7]=1;  end 
14'h 357: begin refPos[0]=43; refFlag[0]=1; refPos[1]=44; refFlag[1]=1; refPos[2]=45; refFlag[2]=1; refPos[3]=46; refFlag[3]=1; refPos[4]=47; refFlag[4]=1; refPos[5]=48; refFlag[5]=1; refPos[6]=49; refFlag[6]=1; refPos[7]=50; refFlag[7]=1;  end 
14'h 360: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=31; refFlag[7]=1;  end 
14'h 361: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=34; refFlag[6]=1; refPos[7]=35; refFlag[7]=1;  end 
14'h 362: begin refPos[0]=31; refFlag[0]=1; refPos[1]=32; refFlag[1]=1; refPos[2]=33; refFlag[2]=1; refPos[3]=34; refFlag[3]=1; refPos[4]=35; refFlag[4]=1; refPos[5]=36; refFlag[5]=1; refPos[6]=37; refFlag[6]=1; refPos[7]=38; refFlag[7]=1;  end 
14'h 363: begin refPos[0]=34; refFlag[0]=1; refPos[1]=35; refFlag[1]=1; refPos[2]=36; refFlag[2]=1; refPos[3]=37; refFlag[3]=1; refPos[4]=38; refFlag[4]=1; refPos[5]=39; refFlag[5]=1; refPos[6]=40; refFlag[6]=1; refPos[7]=41; refFlag[7]=1;  end 
14'h 364: begin refPos[0]=37; refFlag[0]=1; refPos[1]=38; refFlag[1]=1; refPos[2]=39; refFlag[2]=1; refPos[3]=40; refFlag[3]=1; refPos[4]=41; refFlag[4]=1; refPos[5]=42; refFlag[5]=1; refPos[6]=43; refFlag[6]=1; refPos[7]=44; refFlag[7]=1;  end 
14'h 365: begin refPos[0]=41; refFlag[0]=1; refPos[1]=42; refFlag[1]=1; refPos[2]=43; refFlag[2]=1; refPos[3]=44; refFlag[3]=1; refPos[4]=45; refFlag[4]=1; refPos[5]=46; refFlag[5]=1; refPos[6]=47; refFlag[6]=1; refPos[7]=48; refFlag[7]=1;  end 
14'h 366: begin refPos[0]=44; refFlag[0]=1; refPos[1]=45; refFlag[1]=1; refPos[2]=46; refFlag[2]=1; refPos[3]=47; refFlag[3]=1; refPos[4]=48; refFlag[4]=1; refPos[5]=49; refFlag[5]=1; refPos[6]=50; refFlag[6]=1; refPos[7]=51; refFlag[7]=1;  end 
14'h 367: begin refPos[0]=47; refFlag[0]=1; refPos[1]=48; refFlag[1]=1; refPos[2]=49; refFlag[2]=1; refPos[3]=50; refFlag[3]=1; refPos[4]=51; refFlag[4]=1; refPos[5]=52; refFlag[5]=1; refPos[6]=53; refFlag[6]=1; refPos[7]=54; refFlag[7]=1;  end 
14'h 370: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=34; refFlag[6]=1; refPos[7]=35; refFlag[7]=1;  end 
14'h 371: begin refPos[0]=32; refFlag[0]=1; refPos[1]=33; refFlag[1]=1; refPos[2]=34; refFlag[2]=1; refPos[3]=35; refFlag[3]=1; refPos[4]=36; refFlag[4]=1; refPos[5]=37; refFlag[5]=1; refPos[6]=38; refFlag[6]=1; refPos[7]=39; refFlag[7]=1;  end 
14'h 372: begin refPos[0]=35; refFlag[0]=1; refPos[1]=36; refFlag[1]=1; refPos[2]=37; refFlag[2]=1; refPos[3]=38; refFlag[3]=1; refPos[4]=39; refFlag[4]=1; refPos[5]=40; refFlag[5]=1; refPos[6]=41; refFlag[6]=1; refPos[7]=42; refFlag[7]=1;  end 
14'h 373: begin refPos[0]=38; refFlag[0]=1; refPos[1]=39; refFlag[1]=1; refPos[2]=40; refFlag[2]=1; refPos[3]=41; refFlag[3]=1; refPos[4]=42; refFlag[4]=1; refPos[5]=43; refFlag[5]=1; refPos[6]=44; refFlag[6]=1; refPos[7]=45; refFlag[7]=1;  end 
14'h 374: begin refPos[0]=41; refFlag[0]=1; refPos[1]=42; refFlag[1]=1; refPos[2]=43; refFlag[2]=1; refPos[3]=44; refFlag[3]=1; refPos[4]=45; refFlag[4]=1; refPos[5]=46; refFlag[5]=1; refPos[6]=47; refFlag[6]=1; refPos[7]=48; refFlag[7]=1;  end 
14'h 375: begin refPos[0]=45; refFlag[0]=1; refPos[1]=46; refFlag[1]=1; refPos[2]=47; refFlag[2]=1; refPos[3]=48; refFlag[3]=1; refPos[4]=49; refFlag[4]=1; refPos[5]=50; refFlag[5]=1; refPos[6]=51; refFlag[6]=1; refPos[7]=52; refFlag[7]=1;  end 
14'h 376: begin refPos[0]=48; refFlag[0]=1; refPos[1]=49; refFlag[1]=1; refPos[2]=50; refFlag[2]=1; refPos[3]=51; refFlag[3]=1; refPos[4]=52; refFlag[4]=1; refPos[5]=53; refFlag[5]=1; refPos[6]=54; refFlag[6]=1; refPos[7]=55; refFlag[7]=1;  end 
14'h 377: begin refPos[0]=51; refFlag[0]=1; refPos[1]=52; refFlag[1]=1; refPos[2]=53; refFlag[2]=1; refPos[3]=54; refFlag[3]=1; refPos[4]=55; refFlag[4]=1; refPos[5]=56; refFlag[5]=1; refPos[6]=57; refFlag[6]=1; refPos[7]=58; refFlag[7]=1;  end 
14'h 400: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 401: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=9; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 402: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 403: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 404: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 405: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 406: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 407: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=25; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 410: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 411: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=13; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 412: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=15; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 413: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 414: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=21; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 415: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 416: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 417: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=29; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 420: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 421: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 422: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 423: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 424: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=25; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 425: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 426: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 427: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=32; refFlag[5]=1; refPos[6]=33; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 430: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 431: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=21; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 432: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 433: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 434: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=29; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 435: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=31; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 436: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=34; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 437: begin refPos[0]=31; refFlag[0]=1; refPos[1]=32; refFlag[1]=1; refPos[2]=33; refFlag[2]=1; refPos[3]=34; refFlag[3]=1; refPos[4]=35; refFlag[4]=1; refPos[5]=36; refFlag[5]=1; refPos[6]=37; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 440: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 441: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=25; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 442: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 443: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 444: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=32; refFlag[5]=1; refPos[6]=33; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 445: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=35; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 446: begin refPos[0]=32; refFlag[0]=1; refPos[1]=33; refFlag[1]=1; refPos[2]=34; refFlag[2]=1; refPos[3]=35; refFlag[3]=1; refPos[4]=36; refFlag[4]=1; refPos[5]=37; refFlag[5]=1; refPos[6]=38; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 447: begin refPos[0]=35; refFlag[0]=1; refPos[1]=36; refFlag[1]=1; refPos[2]=37; refFlag[2]=1; refPos[3]=38; refFlag[3]=1; refPos[4]=39; refFlag[4]=1; refPos[5]=40; refFlag[5]=1; refPos[6]=41; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 450: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 451: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=29; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 452: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=31; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 453: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=34; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 454: begin refPos[0]=31; refFlag[0]=1; refPos[1]=32; refFlag[1]=1; refPos[2]=33; refFlag[2]=1; refPos[3]=34; refFlag[3]=1; refPos[4]=35; refFlag[4]=1; refPos[5]=36; refFlag[5]=1; refPos[6]=37; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 455: begin refPos[0]=33; refFlag[0]=1; refPos[1]=34; refFlag[1]=1; refPos[2]=35; refFlag[2]=1; refPos[3]=36; refFlag[3]=1; refPos[4]=37; refFlag[4]=1; refPos[5]=38; refFlag[5]=1; refPos[6]=39; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 456: begin refPos[0]=36; refFlag[0]=1; refPos[1]=37; refFlag[1]=1; refPos[2]=38; refFlag[2]=1; refPos[3]=39; refFlag[3]=1; refPos[4]=40; refFlag[4]=1; refPos[5]=41; refFlag[5]=1; refPos[6]=42; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 457: begin refPos[0]=39; refFlag[0]=1; refPos[1]=40; refFlag[1]=1; refPos[2]=41; refFlag[2]=1; refPos[3]=42; refFlag[3]=1; refPos[4]=43; refFlag[4]=1; refPos[5]=44; refFlag[5]=1; refPos[6]=45; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 460: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 461: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=32; refFlag[5]=1; refPos[6]=33; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 462: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=35; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 463: begin refPos[0]=32; refFlag[0]=1; refPos[1]=33; refFlag[1]=1; refPos[2]=34; refFlag[2]=1; refPos[3]=35; refFlag[3]=1; refPos[4]=36; refFlag[4]=1; refPos[5]=37; refFlag[5]=1; refPos[6]=38; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 464: begin refPos[0]=35; refFlag[0]=1; refPos[1]=36; refFlag[1]=1; refPos[2]=37; refFlag[2]=1; refPos[3]=38; refFlag[3]=1; refPos[4]=39; refFlag[4]=1; refPos[5]=40; refFlag[5]=1; refPos[6]=41; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 465: begin refPos[0]=37; refFlag[0]=1; refPos[1]=38; refFlag[1]=1; refPos[2]=39; refFlag[2]=1; refPos[3]=40; refFlag[3]=1; refPos[4]=41; refFlag[4]=1; refPos[5]=42; refFlag[5]=1; refPos[6]=43; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 466: begin refPos[0]=40; refFlag[0]=1; refPos[1]=41; refFlag[1]=1; refPos[2]=42; refFlag[2]=1; refPos[3]=43; refFlag[3]=1; refPos[4]=44; refFlag[4]=1; refPos[5]=45; refFlag[5]=1; refPos[6]=46; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 467: begin refPos[0]=43; refFlag[0]=1; refPos[1]=44; refFlag[1]=1; refPos[2]=45; refFlag[2]=1; refPos[3]=46; refFlag[3]=1; refPos[4]=47; refFlag[4]=1; refPos[5]=48; refFlag[5]=1; refPos[6]=49; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 470: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=34; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 471: begin refPos[0]=31; refFlag[0]=1; refPos[1]=32; refFlag[1]=1; refPos[2]=33; refFlag[2]=1; refPos[3]=34; refFlag[3]=1; refPos[4]=35; refFlag[4]=1; refPos[5]=36; refFlag[5]=1; refPos[6]=37; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 472: begin refPos[0]=33; refFlag[0]=1; refPos[1]=34; refFlag[1]=1; refPos[2]=35; refFlag[2]=1; refPos[3]=36; refFlag[3]=1; refPos[4]=37; refFlag[4]=1; refPos[5]=38; refFlag[5]=1; refPos[6]=39; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 473: begin refPos[0]=36; refFlag[0]=1; refPos[1]=37; refFlag[1]=1; refPos[2]=38; refFlag[2]=1; refPos[3]=39; refFlag[3]=1; refPos[4]=40; refFlag[4]=1; refPos[5]=41; refFlag[5]=1; refPos[6]=42; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 474: begin refPos[0]=39; refFlag[0]=1; refPos[1]=40; refFlag[1]=1; refPos[2]=41; refFlag[2]=1; refPos[3]=42; refFlag[3]=1; refPos[4]=43; refFlag[4]=1; refPos[5]=44; refFlag[5]=1; refPos[6]=45; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 475: begin refPos[0]=41; refFlag[0]=1; refPos[1]=42; refFlag[1]=1; refPos[2]=43; refFlag[2]=1; refPos[3]=44; refFlag[3]=1; refPos[4]=45; refFlag[4]=1; refPos[5]=46; refFlag[5]=1; refPos[6]=47; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 476: begin refPos[0]=44; refFlag[0]=1; refPos[1]=45; refFlag[1]=1; refPos[2]=46; refFlag[2]=1; refPos[3]=47; refFlag[3]=1; refPos[4]=48; refFlag[4]=1; refPos[5]=49; refFlag[5]=1; refPos[6]=50; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 477: begin refPos[0]=47; refFlag[0]=1; refPos[1]=48; refFlag[1]=1; refPos[2]=49; refFlag[2]=1; refPos[3]=50; refFlag[3]=1; refPos[4]=51; refFlag[4]=1; refPos[5]=52; refFlag[5]=1; refPos[6]=53; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 500: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 501: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=8; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 502: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 503: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=12; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 504: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=15; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 505: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 506: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 507: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=21; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 510: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 511: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=12; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 512: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 513: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=16; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 514: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 515: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=21; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 516: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 517: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=25; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 520: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 521: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=16; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 522: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 523: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=20; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 524: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 525: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=25; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 526: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 527: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=29; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 530: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 531: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=20; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 532: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 533: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=24; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 534: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 535: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=29; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 536: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=31; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 537: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=32; refFlag[5]=1; refPos[6]=33; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 540: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 541: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=24; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 542: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 543: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=27; refFlag[5]=1; refPos[6]=28; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 544: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=31; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 545: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=32; refFlag[5]=1; refPos[6]=33; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 546: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=35; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 547: begin refPos[0]=31; refFlag[0]=1; refPos[1]=32; refFlag[1]=1; refPos[2]=33; refFlag[2]=1; refPos[3]=34; refFlag[3]=1; refPos[4]=35; refFlag[4]=1; refPos[5]=36; refFlag[5]=1; refPos[6]=37; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 550: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 551: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=27; refFlag[5]=1; refPos[6]=28; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 552: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 553: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=31; refFlag[5]=1; refPos[6]=32; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 554: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=35; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 555: begin refPos[0]=31; refFlag[0]=1; refPos[1]=32; refFlag[1]=1; refPos[2]=33; refFlag[2]=1; refPos[3]=34; refFlag[3]=1; refPos[4]=35; refFlag[4]=1; refPos[5]=36; refFlag[5]=1; refPos[6]=37; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 556: begin refPos[0]=33; refFlag[0]=1; refPos[1]=34; refFlag[1]=1; refPos[2]=35; refFlag[2]=1; refPos[3]=36; refFlag[3]=1; refPos[4]=37; refFlag[4]=1; refPos[5]=38; refFlag[5]=1; refPos[6]=39; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 557: begin refPos[0]=35; refFlag[0]=1; refPos[1]=36; refFlag[1]=1; refPos[2]=37; refFlag[2]=1; refPos[3]=38; refFlag[3]=1; refPos[4]=39; refFlag[4]=1; refPos[5]=40; refFlag[5]=1; refPos[6]=41; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 560: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 561: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=31; refFlag[5]=1; refPos[6]=32; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 562: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=34; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 563: begin refPos[0]=30; refFlag[0]=1; refPos[1]=31; refFlag[1]=1; refPos[2]=32; refFlag[2]=1; refPos[3]=33; refFlag[3]=1; refPos[4]=34; refFlag[4]=1; refPos[5]=35; refFlag[5]=1; refPos[6]=36; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 564: begin refPos[0]=33; refFlag[0]=1; refPos[1]=34; refFlag[1]=1; refPos[2]=35; refFlag[2]=1; refPos[3]=36; refFlag[3]=1; refPos[4]=37; refFlag[4]=1; refPos[5]=38; refFlag[5]=1; refPos[6]=39; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 565: begin refPos[0]=35; refFlag[0]=1; refPos[1]=36; refFlag[1]=1; refPos[2]=37; refFlag[2]=1; refPos[3]=38; refFlag[3]=1; refPos[4]=39; refFlag[4]=1; refPos[5]=40; refFlag[5]=1; refPos[6]=41; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 566: begin refPos[0]=37; refFlag[0]=1; refPos[1]=38; refFlag[1]=1; refPos[2]=39; refFlag[2]=1; refPos[3]=40; refFlag[3]=1; refPos[4]=41; refFlag[4]=1; refPos[5]=42; refFlag[5]=1; refPos[6]=43; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 567: begin refPos[0]=39; refFlag[0]=1; refPos[1]=40; refFlag[1]=1; refPos[2]=41; refFlag[2]=1; refPos[3]=42; refFlag[3]=1; refPos[4]=43; refFlag[4]=1; refPos[5]=44; refFlag[5]=1; refPos[6]=45; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 570: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=34; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 571: begin refPos[0]=30; refFlag[0]=1; refPos[1]=31; refFlag[1]=1; refPos[2]=32; refFlag[2]=1; refPos[3]=33; refFlag[3]=1; refPos[4]=34; refFlag[4]=1; refPos[5]=35; refFlag[5]=1; refPos[6]=36; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 572: begin refPos[0]=32; refFlag[0]=1; refPos[1]=33; refFlag[1]=1; refPos[2]=34; refFlag[2]=1; refPos[3]=35; refFlag[3]=1; refPos[4]=36; refFlag[4]=1; refPos[5]=37; refFlag[5]=1; refPos[6]=38; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 573: begin refPos[0]=34; refFlag[0]=1; refPos[1]=35; refFlag[1]=1; refPos[2]=36; refFlag[2]=1; refPos[3]=37; refFlag[3]=1; refPos[4]=38; refFlag[4]=1; refPos[5]=39; refFlag[5]=1; refPos[6]=40; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 574: begin refPos[0]=37; refFlag[0]=1; refPos[1]=38; refFlag[1]=1; refPos[2]=39; refFlag[2]=1; refPos[3]=40; refFlag[3]=1; refPos[4]=41; refFlag[4]=1; refPos[5]=42; refFlag[5]=1; refPos[6]=43; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 575: begin refPos[0]=39; refFlag[0]=1; refPos[1]=40; refFlag[1]=1; refPos[2]=41; refFlag[2]=1; refPos[3]=42; refFlag[3]=1; refPos[4]=43; refFlag[4]=1; refPos[5]=44; refFlag[5]=1; refPos[6]=45; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 576: begin refPos[0]=41; refFlag[0]=1; refPos[1]=42; refFlag[1]=1; refPos[2]=43; refFlag[2]=1; refPos[3]=44; refFlag[3]=1; refPos[4]=45; refFlag[4]=1; refPos[5]=46; refFlag[5]=1; refPos[6]=47; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 577: begin refPos[0]=43; refFlag[0]=1; refPos[1]=44; refFlag[1]=1; refPos[2]=45; refFlag[2]=1; refPos[3]=46; refFlag[3]=1; refPos[4]=47; refFlag[4]=1; refPos[5]=48; refFlag[5]=1; refPos[6]=49; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 600: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 601: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=8; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 602: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=9; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 603: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 604: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=12; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 605: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 606: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=16; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 607: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 610: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 611: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=12; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 612: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=13; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 613: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=15; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 614: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=16; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 615: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 616: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=20; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 617: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=21; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 620: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 621: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=16; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 622: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 623: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 624: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=20; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 625: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 626: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=24; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 627: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=25; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 630: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 631: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=20; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 632: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=21; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 633: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 634: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=24; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 635: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 636: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=27; refFlag[5]=1; refPos[6]=28; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 637: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=29; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 640: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 641: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=24; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 642: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=25; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 643: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 644: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=27; refFlag[5]=1; refPos[6]=28; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 645: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 646: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=31; refFlag[5]=1; refPos[6]=32; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 647: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=32; refFlag[5]=1; refPos[6]=33; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 650: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 651: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=27; refFlag[5]=1; refPos[6]=28; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 652: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=29; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 653: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=31; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 654: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=31; refFlag[5]=1; refPos[6]=32; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 655: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=34; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 656: begin refPos[0]=30; refFlag[0]=1; refPos[1]=31; refFlag[1]=1; refPos[2]=32; refFlag[2]=1; refPos[3]=33; refFlag[3]=1; refPos[4]=34; refFlag[4]=1; refPos[5]=35; refFlag[5]=1; refPos[6]=36; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 657: begin refPos[0]=31; refFlag[0]=1; refPos[1]=32; refFlag[1]=1; refPos[2]=33; refFlag[2]=1; refPos[3]=34; refFlag[3]=1; refPos[4]=35; refFlag[4]=1; refPos[5]=36; refFlag[5]=1; refPos[6]=37; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 660: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 661: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=31; refFlag[5]=1; refPos[6]=32; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 662: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=32; refFlag[5]=1; refPos[6]=33; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 663: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=35; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 664: begin refPos[0]=30; refFlag[0]=1; refPos[1]=31; refFlag[1]=1; refPos[2]=32; refFlag[2]=1; refPos[3]=33; refFlag[3]=1; refPos[4]=34; refFlag[4]=1; refPos[5]=35; refFlag[5]=1; refPos[6]=36; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 665: begin refPos[0]=32; refFlag[0]=1; refPos[1]=33; refFlag[1]=1; refPos[2]=34; refFlag[2]=1; refPos[3]=35; refFlag[3]=1; refPos[4]=36; refFlag[4]=1; refPos[5]=37; refFlag[5]=1; refPos[6]=38; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 666: begin refPos[0]=34; refFlag[0]=1; refPos[1]=35; refFlag[1]=1; refPos[2]=36; refFlag[2]=1; refPos[3]=37; refFlag[3]=1; refPos[4]=38; refFlag[4]=1; refPos[5]=39; refFlag[5]=1; refPos[6]=40; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 667: begin refPos[0]=35; refFlag[0]=1; refPos[1]=36; refFlag[1]=1; refPos[2]=37; refFlag[2]=1; refPos[3]=38; refFlag[3]=1; refPos[4]=39; refFlag[4]=1; refPos[5]=40; refFlag[5]=1; refPos[6]=41; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 670: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=34; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 671: begin refPos[0]=30; refFlag[0]=1; refPos[1]=31; refFlag[1]=1; refPos[2]=32; refFlag[2]=1; refPos[3]=33; refFlag[3]=1; refPos[4]=34; refFlag[4]=1; refPos[5]=35; refFlag[5]=1; refPos[6]=36; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 672: begin refPos[0]=31; refFlag[0]=1; refPos[1]=32; refFlag[1]=1; refPos[2]=33; refFlag[2]=1; refPos[3]=34; refFlag[3]=1; refPos[4]=35; refFlag[4]=1; refPos[5]=36; refFlag[5]=1; refPos[6]=37; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 673: begin refPos[0]=33; refFlag[0]=1; refPos[1]=34; refFlag[1]=1; refPos[2]=35; refFlag[2]=1; refPos[3]=36; refFlag[3]=1; refPos[4]=37; refFlag[4]=1; refPos[5]=38; refFlag[5]=1; refPos[6]=39; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 674: begin refPos[0]=34; refFlag[0]=1; refPos[1]=35; refFlag[1]=1; refPos[2]=36; refFlag[2]=1; refPos[3]=37; refFlag[3]=1; refPos[4]=38; refFlag[4]=1; refPos[5]=39; refFlag[5]=1; refPos[6]=40; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 675: begin refPos[0]=36; refFlag[0]=1; refPos[1]=37; refFlag[1]=1; refPos[2]=38; refFlag[2]=1; refPos[3]=39; refFlag[3]=1; refPos[4]=40; refFlag[4]=1; refPos[5]=41; refFlag[5]=1; refPos[6]=42; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 676: begin refPos[0]=38; refFlag[0]=1; refPos[1]=39; refFlag[1]=1; refPos[2]=40; refFlag[2]=1; refPos[3]=41; refFlag[3]=1; refPos[4]=42; refFlag[4]=1; refPos[5]=43; refFlag[5]=1; refPos[6]=44; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 677: begin refPos[0]=39; refFlag[0]=1; refPos[1]=40; refFlag[1]=1; refPos[2]=41; refFlag[2]=1; refPos[3]=42; refFlag[3]=1; refPos[4]=43; refFlag[4]=1; refPos[5]=44; refFlag[5]=1; refPos[6]=45; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 700: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 701: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 702: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 703: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 704: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 705: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 706: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 707: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 710: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 711: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 712: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 713: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 714: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 715: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 716: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 717: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 720: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 721: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 722: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 723: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 724: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 725: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 726: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 727: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 730: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 731: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 732: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 733: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 734: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 735: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 736: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 737: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 740: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 741: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 742: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 743: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 744: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 745: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 746: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 747: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 750: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 751: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 752: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=27; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 753: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 754: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 755: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 756: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=32; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 757: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 760: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 761: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 762: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=31; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 763: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=32; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 764: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 765: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 766: begin refPos[0]=31; refFlag[0]=1; refPos[1]=32; refFlag[1]=1; refPos[2]=33; refFlag[2]=1; refPos[3]=34; refFlag[3]=1; refPos[4]=35; refFlag[4]=1; refPos[5]=36; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 767: begin refPos[0]=32; refFlag[0]=1; refPos[1]=33; refFlag[1]=1; refPos[2]=34; refFlag[2]=1; refPos[3]=35; refFlag[3]=1; refPos[4]=36; refFlag[4]=1; refPos[5]=37; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 770: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 771: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 772: begin refPos[0]=30; refFlag[0]=1; refPos[1]=31; refFlag[1]=1; refPos[2]=32; refFlag[2]=1; refPos[3]=33; refFlag[3]=1; refPos[4]=34; refFlag[4]=1; refPos[5]=35; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 773: begin refPos[0]=31; refFlag[0]=1; refPos[1]=32; refFlag[1]=1; refPos[2]=33; refFlag[2]=1; refPos[3]=34; refFlag[3]=1; refPos[4]=35; refFlag[4]=1; refPos[5]=36; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 774: begin refPos[0]=32; refFlag[0]=1; refPos[1]=33; refFlag[1]=1; refPos[2]=34; refFlag[2]=1; refPos[3]=35; refFlag[3]=1; refPos[4]=36; refFlag[4]=1; refPos[5]=37; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 775: begin refPos[0]=33; refFlag[0]=1; refPos[1]=34; refFlag[1]=1; refPos[2]=35; refFlag[2]=1; refPos[3]=36; refFlag[3]=1; refPos[4]=37; refFlag[4]=1; refPos[5]=38; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 776: begin refPos[0]=35; refFlag[0]=1; refPos[1]=36; refFlag[1]=1; refPos[2]=37; refFlag[2]=1; refPos[3]=38; refFlag[3]=1; refPos[4]=39; refFlag[4]=1; refPos[5]=40; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 777: begin refPos[0]=36; refFlag[0]=1; refPos[1]=37; refFlag[1]=1; refPos[2]=38; refFlag[2]=1; refPos[3]=39; refFlag[3]=1; refPos[4]=40; refFlag[4]=1; refPos[5]=41; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 800: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 801: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 802: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 803: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 804: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 805: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 806: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 807: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 810: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 811: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 812: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 813: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 814: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 815: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 816: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 817: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 820: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 821: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 822: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 823: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 824: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 825: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 826: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 827: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 830: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 831: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 832: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 833: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 834: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 835: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 836: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 837: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 840: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 841: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 842: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 843: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 844: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 845: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 846: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 847: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 850: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 851: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 852: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 853: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=27; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 854: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=27; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 855: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 856: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 857: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 860: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 861: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 862: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 863: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=31; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 864: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=31; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 865: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=32; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 866: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=32; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 867: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 870: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 871: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 872: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 873: begin refPos[0]=30; refFlag[0]=1; refPos[1]=31; refFlag[1]=1; refPos[2]=32; refFlag[2]=1; refPos[3]=33; refFlag[3]=1; refPos[4]=34; refFlag[4]=1; refPos[5]=35; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 874: begin refPos[0]=30; refFlag[0]=1; refPos[1]=31; refFlag[1]=1; refPos[2]=32; refFlag[2]=1; refPos[3]=33; refFlag[3]=1; refPos[4]=34; refFlag[4]=1; refPos[5]=35; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 875: begin refPos[0]=31; refFlag[0]=1; refPos[1]=32; refFlag[1]=1; refPos[2]=33; refFlag[2]=1; refPos[3]=34; refFlag[3]=1; refPos[4]=35; refFlag[4]=1; refPos[5]=36; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 876: begin refPos[0]=31; refFlag[0]=1; refPos[1]=32; refFlag[1]=1; refPos[2]=33; refFlag[2]=1; refPos[3]=34; refFlag[3]=1; refPos[4]=35; refFlag[4]=1; refPos[5]=36; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 877: begin refPos[0]=32; refFlag[0]=1; refPos[1]=33; refFlag[1]=1; refPos[2]=34; refFlag[2]=1; refPos[3]=35; refFlag[3]=1; refPos[4]=36; refFlag[4]=1; refPos[5]=37; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 900: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 901: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 902: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 903: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 904: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 905: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 906: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 907: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 910: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 911: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 912: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 913: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 914: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 915: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 916: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 917: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 920: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 921: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 922: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 923: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 924: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 925: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 926: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 927: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 930: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 931: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 932: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 933: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 934: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 935: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 936: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 937: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 940: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 941: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 942: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 943: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 944: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 945: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 946: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 947: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 950: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 951: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 952: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 953: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 954: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 955: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 956: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 957: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 960: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 961: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 962: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 963: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 964: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 965: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 966: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 967: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 970: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 971: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 972: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 973: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=32; refFlag[4]=1; refPos[5]=33; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 974: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 975: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 976: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h 977: begin refPos[0]=29; refFlag[0]=1; refPos[1]=30; refFlag[1]=1; refPos[2]=31; refFlag[2]=1; refPos[3]=32; refFlag[3]=1; refPos[4]=33; refFlag[4]=1; refPos[5]=34; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a00: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=2; refFlag[6]=0; refPos[7]=3; refFlag[7]=0;  end 
14'h a01: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=7; refFlag[7]=0;  end 
14'h a02: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=11; refFlag[7]=0;  end 
14'h a03: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=15; refFlag[7]=0;  end 
14'h a04: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a05: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a06: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a07: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a10: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a11: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a12: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a13: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a14: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a15: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a16: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a17: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a20: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a21: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a22: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a23: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a24: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a25: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a26: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a27: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a30: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a31: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a32: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a33: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a34: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a35: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a36: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a37: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a40: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a41: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a42: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a43: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a44: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a45: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a46: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a47: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a50: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a51: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a52: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a53: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a54: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a55: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a56: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a57: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a60: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a61: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a62: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a63: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a64: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a65: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a66: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a67: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a70: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a71: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a72: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a73: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a74: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a75: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a76: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h a77: begin refPos[0]=28; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=30; refFlag[2]=1; refPos[3]=31; refFlag[3]=1; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b00: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b01: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b02: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b03: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b04: begin refPos[0]=15; refFlag[0]=0; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b05: begin refPos[0]=15; refFlag[0]=0; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b06: begin refPos[0]=15; refFlag[0]=0; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b07: begin refPos[0]=15; refFlag[0]=0; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b10: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b11: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b12: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b13: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b14: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b15: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b16: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b17: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b20: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b21: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b22: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b23: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b24: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b25: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b26: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b27: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b30: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b31: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b32: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b33: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b34: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b35: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b36: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b37: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b40: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b41: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b42: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b43: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b44: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b45: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b46: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b47: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b50: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b51: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b52: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b53: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b54: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b55: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b56: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b57: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b60: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b61: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b62: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b63: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b64: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b65: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b66: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b67: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b70: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b71: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b72: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b73: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b74: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b75: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b76: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h b77: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c00: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c01: begin refPos[0]=5; refFlag[0]=0; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=3; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c02: begin refPos[0]=5; refFlag[0]=0; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=3; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c03: begin refPos[0]=12; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=2; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c04: begin refPos[0]=18; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c05: begin refPos[0]=18; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c06: begin refPos[0]=25; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c07: begin refPos[0]=25; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c10: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c11: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c12: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c13: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c14: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c15: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c16: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c17: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c20: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c21: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c22: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c23: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c24: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c25: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c26: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c27: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c30: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c31: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c32: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c33: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c34: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c35: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c36: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c37: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c40: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c41: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c42: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c43: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c44: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c45: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c46: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c47: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c50: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c51: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c52: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c53: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c54: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c55: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c56: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c57: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c60: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c61: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=27; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c62: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=27; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c63: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c64: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c65: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c66: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c67: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c70: begin refPos[0]=27; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=29; refFlag[2]=1; refPos[3]=30; refFlag[3]=1; refPos[4]=31; refFlag[4]=1; refPos[5]=32; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c71: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=31; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c72: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=31; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c73: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c74: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c75: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c76: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h c77: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d00: begin refPos[0]=3; refFlag[0]=0; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=3; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d01: begin refPos[0]=6; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=2; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d02: begin refPos[0]=10; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d03: begin refPos[0]=13; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d04: begin refPos[0]=17; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=99; refFlag[5]=2; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d05: begin refPos[0]=20; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=3; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d06: begin refPos[0]=24; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d07: begin refPos[0]=27; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d10: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d11: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d12: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d13: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d14: begin refPos[0]=3; refFlag[0]=0; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=3; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d15: begin refPos[0]=6; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=2; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d16: begin refPos[0]=10; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d17: begin refPos[0]=13; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d20: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d21: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d22: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d23: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d24: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d25: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d26: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d27: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d30: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d31: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d32: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d33: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d34: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d35: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d36: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d37: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d40: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d41: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d42: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d43: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d44: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d45: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d46: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d47: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d50: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d51: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d52: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d53: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d54: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d55: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d56: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d57: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d60: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=27; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d61: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d62: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d63: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d64: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d65: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d66: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d67: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d70: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=31; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d71: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d72: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d73: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d74: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=27; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d75: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d76: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h d77: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e00: begin refPos[0]=1; refFlag[0]=0; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=3; refFlag[5]=1; refPos[6]=4; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e01: begin refPos[0]=6; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e02: begin refPos[0]=9; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=1; refPos[6]=1; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e03: begin refPos[0]=14; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=99; refFlag[6]=2; refPos[7]=1; refFlag[7]=-1;  end 
14'h e04: begin refPos[0]=19; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=4; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h e05: begin refPos[0]=21; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h e06: begin refPos[0]=26; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h e07: begin refPos[0]=29; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h e10: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=8; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e11: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e12: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=5; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e13: begin refPos[0]=4; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=2; refFlag[5]=1; refPos[6]=3; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e14: begin refPos[0]=9; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=1; refPos[6]=1; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e15: begin refPos[0]=11; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=99; refFlag[5]=2; refPos[6]=0; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e16: begin refPos[0]=16; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h e17: begin refPos[0]=19; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=4; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h e20: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=12; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e21: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e22: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=9; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e23: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=7; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e24: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=5; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e25: begin refPos[0]=1; refFlag[0]=0; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=3; refFlag[5]=1; refPos[6]=4; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e26: begin refPos[0]=6; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e27: begin refPos[0]=9; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=1; refPos[6]=1; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e30: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=16; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e31: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e32: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=13; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e33: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e34: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=9; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e35: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=8; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e36: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e37: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=5; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e40: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=20; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e41: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e42: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e43: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=15; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e44: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=13; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e45: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=12; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e46: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e47: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=9; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e50: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=24; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e51: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e52: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=21; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e53: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e54: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e55: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=16; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e56: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e57: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=13; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e60: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=27; refFlag[5]=1; refPos[6]=28; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e61: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e62: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=25; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e63: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e64: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=21; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e65: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=20; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e66: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e67: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e70: begin refPos[0]=26; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=29; refFlag[3]=1; refPos[4]=30; refFlag[4]=1; refPos[5]=31; refFlag[5]=1; refPos[6]=32; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e71: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e72: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=29; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e73: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e74: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=25; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e75: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=24; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e76: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h e77: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=21; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f00: begin refPos[0]=3; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=2; refFlag[5]=1; refPos[6]=3; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f01: begin refPos[0]=7; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=1; refPos[6]=1; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f02: begin refPos[0]=10; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=99; refFlag[6]=2; refPos[7]=1; refFlag[7]=-1;  end 
14'h f03: begin refPos[0]=14; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=3; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h f04: begin refPos[0]=18; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=7; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h f05: begin refPos[0]=22; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h f06: begin refPos[0]=25; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h f07: begin refPos[0]=29; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h f10: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=7; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f11: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=5; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f12: begin refPos[0]=3; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=2; refFlag[5]=1; refPos[6]=3; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f13: begin refPos[0]=7; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=1; refPos[6]=1; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f14: begin refPos[0]=10; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=99; refFlag[6]=2; refPos[7]=1; refFlag[7]=-1;  end 
14'h f15: begin refPos[0]=14; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=3; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h f16: begin refPos[0]=18; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=7; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h f17: begin refPos[0]=22; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h f20: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f21: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=9; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f22: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=7; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f23: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=5; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f24: begin refPos[0]=3; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=2; refFlag[5]=1; refPos[6]=3; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f25: begin refPos[0]=7; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=1; refPos[6]=1; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f26: begin refPos[0]=10; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=99; refFlag[6]=2; refPos[7]=1; refFlag[7]=-1;  end 
14'h f27: begin refPos[0]=14; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=3; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h f30: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=15; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f31: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=13; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f32: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f33: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=9; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f34: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=7; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f35: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=5; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f36: begin refPos[0]=3; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=2; refFlag[5]=1; refPos[6]=3; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f37: begin refPos[0]=7; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=1; refPos[6]=1; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f40: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f41: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f42: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=15; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f43: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=13; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f44: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f45: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=9; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f46: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=7; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f47: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=5; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f50: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f51: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=21; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f52: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f53: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f54: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=15; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f55: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=13; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f56: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f57: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=9; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f60: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f61: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=25; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f62: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f63: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=21; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f64: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f65: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f66: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=15; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f67: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=13; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f70: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=31; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f71: begin refPos[0]=23; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=27; refFlag[4]=1; refPos[5]=28; refFlag[5]=1; refPos[6]=29; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f72: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f73: begin refPos[0]=19; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=25; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f74: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f75: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=21; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f76: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h f77: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1000: begin refPos[0]=2; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=2; refFlag[5]=1; refPos[6]=3; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1001: begin refPos[0]=7; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=99; refFlag[5]=2; refPos[6]=0; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1002: begin refPos[0]=10; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=2; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1003: begin refPos[0]=14; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=5; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1004: begin refPos[0]=19; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1005: begin refPos[0]=22; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=13; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1006: begin refPos[0]=26; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1007: begin refPos[0]=29; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=20; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1010: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=7; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1011: begin refPos[0]=1; refFlag[0]=0; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=3; refFlag[5]=1; refPos[6]=4; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1012: begin refPos[0]=4; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1013: begin refPos[0]=8; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=2; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=99; refFlag[6]=2; refPos[7]=1; refFlag[7]=-1;  end 
14'h1014: begin refPos[0]=13; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=4; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1015: begin refPos[0]=16; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=7; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1016: begin refPos[0]=20; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1017: begin refPos[0]=23; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1020: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1021: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=8; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1022: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1023: begin refPos[0]=2; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=2; refFlag[5]=1; refPos[6]=3; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1024: begin refPos[0]=7; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=99; refFlag[5]=2; refPos[6]=0; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1025: begin refPos[0]=10; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=2; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1026: begin refPos[0]=14; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=5; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1027: begin refPos[0]=17; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=8; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1030: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=15; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1031: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=12; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1032: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1033: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=7; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1034: begin refPos[0]=1; refFlag[0]=0; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=3; refFlag[5]=1; refPos[6]=4; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1035: begin refPos[0]=4; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1036: begin refPos[0]=8; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=2; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=99; refFlag[6]=2; refPos[7]=1; refFlag[7]=-1;  end 
14'h1037: begin refPos[0]=11; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=2; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1040: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1041: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=16; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1042: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1043: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1044: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=8; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1045: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1046: begin refPos[0]=2; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=2; refFlag[5]=1; refPos[6]=3; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1047: begin refPos[0]=5; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=1; refPos[6]=1; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1050: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1051: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=20; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1052: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1053: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=15; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1054: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=12; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1055: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1056: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=7; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1057: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=5; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1060: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1061: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=24; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1062: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1063: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1064: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=16; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1065: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1066: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1067: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=9; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1070: begin refPos[0]=25; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=28; refFlag[3]=1; refPos[4]=29; refFlag[4]=1; refPos[5]=30; refFlag[5]=1; refPos[6]=31; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1071: begin refPos[0]=22; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=27; refFlag[5]=1; refPos[6]=28; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1072: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1073: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1074: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=20; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1075: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1076: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=15; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1077: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=13; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1100: begin refPos[0]=3; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=0; refFlag[2]=0; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h1101: begin refPos[0]=6; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=0; refFlag[5]=0; refPos[6]=99; refFlag[6]=2; refPos[7]=0; refFlag[7]=1;  end 
14'h1102: begin refPos[0]=10; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=3; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h1103: begin refPos[0]=14; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=5; refFlag[7]=0;  end 
14'h1104: begin refPos[0]=19; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=10; refFlag[7]=0;  end 
14'h1105: begin refPos[0]=22; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=15; refFlag[6]=0; refPos[7]=14; refFlag[7]=0;  end 
14'h1106: begin refPos[0]=26; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=17; refFlag[7]=0;  end 
14'h1107: begin refPos[0]=30; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=21; refFlag[7]=0;  end 
14'h1110: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h1111: begin refPos[0]=1; refFlag[0]=0; refPos[1]=0; refFlag[1]=0; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=2; refFlag[5]=1; refPos[6]=3; refFlag[6]=1; refPos[7]=4; refFlag[7]=1;  end 
14'h1112: begin refPos[0]=5; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=0; refFlag[4]=0; refPos[5]=99; refFlag[5]=2; refPos[6]=0; refFlag[6]=1; refPos[7]=1; refFlag[7]=1;  end 
14'h1113: begin refPos[0]=9; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=3; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=0; refFlag[7]=0;  end 
14'h1114: begin refPos[0]=14; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=5; refFlag[7]=0;  end 
14'h1115: begin refPos[0]=17; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=9; refFlag[7]=0;  end 
14'h1116: begin refPos[0]=21; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=13; refFlag[7]=0;  end 
14'h1117: begin refPos[0]=25; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=16; refFlag[7]=0;  end 
14'h1120: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h1121: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=7; refFlag[6]=1; refPos[7]=8; refFlag[7]=1;  end 
14'h1122: begin refPos[0]=0; refFlag[0]=0; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=3; refFlag[5]=1; refPos[6]=4; refFlag[6]=1; refPos[7]=5; refFlag[7]=1;  end 
14'h1123: begin refPos[0]=4; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=0; refFlag[3]=0; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=1; refPos[6]=1; refFlag[6]=1; refPos[7]=2; refFlag[7]=1;  end 
14'h1124: begin refPos[0]=9; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=3; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=0; refFlag[7]=0;  end 
14'h1125: begin refPos[0]=13; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=5; refFlag[6]=0; refPos[7]=4; refFlag[7]=0;  end 
14'h1126: begin refPos[0]=16; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=9; refFlag[6]=0; refPos[7]=8; refFlag[7]=0;  end 
14'h1127: begin refPos[0]=20; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=13; refFlag[6]=0; refPos[7]=11; refFlag[7]=0;  end 
14'h1130: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
14'h1131: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=12; refFlag[7]=1;  end 
14'h1132: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=8; refFlag[6]=1; refPos[7]=9; refFlag[7]=1;  end 
14'h1133: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=5; refFlag[6]=1; refPos[7]=6; refFlag[7]=1;  end 
14'h1134: begin refPos[0]=4; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=0; refFlag[3]=0; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=1; refPos[6]=1; refFlag[6]=1; refPos[7]=2; refFlag[7]=1;  end 
14'h1135: begin refPos[0]=8; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=0; refFlag[6]=0; refPos[7]=99; refFlag[7]=2;  end 
14'h1136: begin refPos[0]=11; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=4; refFlag[6]=0; refPos[7]=3; refFlag[7]=0;  end 
14'h1137: begin refPos[0]=15; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=8; refFlag[6]=0; refPos[7]=6; refFlag[7]=0;  end 
14'h1140: begin refPos[0]=12; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=19; refFlag[7]=1;  end 
14'h1141: begin refPos[0]=9; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=15; refFlag[6]=1; refPos[7]=16; refFlag[7]=1;  end 
14'h1142: begin refPos[0]=6; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=12; refFlag[6]=1; refPos[7]=13; refFlag[7]=1;  end 
14'h1143: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=9; refFlag[6]=1; refPos[7]=10; refFlag[7]=1;  end 
14'h1144: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=5; refFlag[6]=1; refPos[7]=6; refFlag[7]=1;  end 
14'h1145: begin refPos[0]=3; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=0; refFlag[2]=0; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h1146: begin refPos[0]=6; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=0; refFlag[5]=0; refPos[6]=99; refFlag[6]=2; refPos[7]=0; refFlag[7]=1;  end 
14'h1147: begin refPos[0]=10; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=3; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h1150: begin refPos[0]=16; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=23; refFlag[7]=1;  end 
14'h1151: begin refPos[0]=13; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=18; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=20; refFlag[7]=1;  end 
14'h1152: begin refPos[0]=10; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=16; refFlag[6]=1; refPos[7]=17; refFlag[7]=1;  end 
14'h1153: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=13; refFlag[6]=1; refPos[7]=14; refFlag[7]=1;  end 
14'h1154: begin refPos[0]=3; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=9; refFlag[6]=1; refPos[7]=10; refFlag[7]=1;  end 
14'h1155: begin refPos[0]=0; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h1156: begin refPos[0]=1; refFlag[0]=0; refPos[1]=0; refFlag[1]=0; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=2; refFlag[5]=1; refPos[6]=3; refFlag[6]=1; refPos[7]=4; refFlag[7]=1;  end 
14'h1157: begin refPos[0]=5; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=0; refFlag[4]=0; refPos[5]=99; refFlag[5]=2; refPos[6]=0; refFlag[6]=1; refPos[7]=1; refFlag[7]=1;  end 
14'h1160: begin refPos[0]=20; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=24; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=26; refFlag[6]=1; refPos[7]=27; refFlag[7]=1;  end 
14'h1161: begin refPos[0]=17; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=23; refFlag[6]=1; refPos[7]=24; refFlag[7]=1;  end 
14'h1162: begin refPos[0]=14; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=20; refFlag[6]=1; refPos[7]=21; refFlag[7]=1;  end 
14'h1163: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=18; refFlag[7]=1;  end 
14'h1164: begin refPos[0]=7; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=13; refFlag[6]=1; refPos[7]=14; refFlag[7]=1;  end 
14'h1165: begin refPos[0]=4; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h1166: begin refPos[0]=1; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=7; refFlag[6]=1; refPos[7]=8; refFlag[7]=1;  end 
14'h1167: begin refPos[0]=0; refFlag[0]=0; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=3; refFlag[5]=1; refPos[6]=4; refFlag[6]=1; refPos[7]=5; refFlag[7]=1;  end 
14'h1170: begin refPos[0]=24; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=28; refFlag[4]=1; refPos[5]=29; refFlag[5]=1; refPos[6]=30; refFlag[6]=1; refPos[7]=31; refFlag[7]=1;  end 
14'h1171: begin refPos[0]=21; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=24; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=26; refFlag[5]=1; refPos[6]=27; refFlag[6]=1; refPos[7]=28; refFlag[7]=1;  end 
14'h1172: begin refPos[0]=18; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=23; refFlag[5]=1; refPos[6]=24; refFlag[6]=1; refPos[7]=25; refFlag[7]=1;  end 
14'h1173: begin refPos[0]=15; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=18; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=21; refFlag[6]=1; refPos[7]=22; refFlag[7]=1;  end 
14'h1174: begin refPos[0]=11; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=18; refFlag[7]=1;  end 
14'h1175: begin refPos[0]=8; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
14'h1176: begin refPos[0]=5; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=12; refFlag[7]=1;  end 
14'h1177: begin refPos[0]=2; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=8; refFlag[6]=1; refPos[7]=9; refFlag[7]=1;  end 
14'h1200: begin refPos[0]=2; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=0; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=2; refFlag[6]=0; refPos[7]=3; refFlag[7]=0;  end 
14'h1201: begin refPos[0]=6; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=0; refFlag[6]=1; refPos[7]=99; refFlag[7]=2;  end 
14'h1202: begin refPos[0]=10; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=4; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h1203: begin refPos[0]=14; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=8; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h1204: begin refPos[0]=18; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=12; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h1205: begin refPos[0]=22; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=16; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
14'h1206: begin refPos[0]=26; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=20; refFlag[6]=1; refPos[7]=19; refFlag[7]=1;  end 
14'h1207: begin refPos[0]=30; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=28; refFlag[2]=1; refPos[3]=27; refFlag[3]=1; refPos[4]=26; refFlag[4]=1; refPos[5]=25; refFlag[5]=1; refPos[6]=24; refFlag[6]=1; refPos[7]=23; refFlag[7]=1;  end 
14'h1210: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=7; refFlag[7]=0;  end 
14'h1211: begin refPos[0]=2; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=0; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=2; refFlag[6]=0; refPos[7]=3; refFlag[7]=0;  end 
14'h1212: begin refPos[0]=6; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=0; refFlag[6]=1; refPos[7]=99; refFlag[7]=2;  end 
14'h1213: begin refPos[0]=10; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=4; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h1214: begin refPos[0]=14; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=8; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h1215: begin refPos[0]=18; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=12; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h1216: begin refPos[0]=22; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=16; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
14'h1217: begin refPos[0]=26; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=21; refFlag[5]=1; refPos[6]=20; refFlag[6]=1; refPos[7]=19; refFlag[7]=1;  end 
14'h1220: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=11; refFlag[7]=0;  end 
14'h1221: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=7; refFlag[7]=0;  end 
14'h1222: begin refPos[0]=2; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=0; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=2; refFlag[6]=0; refPos[7]=3; refFlag[7]=0;  end 
14'h1223: begin refPos[0]=6; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=0; refFlag[6]=1; refPos[7]=99; refFlag[7]=2;  end 
14'h1224: begin refPos[0]=10; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=4; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h1225: begin refPos[0]=14; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=8; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h1226: begin refPos[0]=18; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=12; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h1227: begin refPos[0]=22; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=17; refFlag[5]=1; refPos[6]=16; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
14'h1230: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=15; refFlag[7]=0;  end 
14'h1231: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=11; refFlag[7]=0;  end 
14'h1232: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=7; refFlag[7]=0;  end 
14'h1233: begin refPos[0]=2; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=0; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=2; refFlag[6]=0; refPos[7]=3; refFlag[7]=0;  end 
14'h1234: begin refPos[0]=6; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=0; refFlag[6]=1; refPos[7]=99; refFlag[7]=2;  end 
14'h1235: begin refPos[0]=10; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=4; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h1236: begin refPos[0]=14; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=8; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h1237: begin refPos[0]=18; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=12; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h1240: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=19; refFlag[7]=0;  end 
14'h1241: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=15; refFlag[7]=0;  end 
14'h1242: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=11; refFlag[7]=0;  end 
14'h1243: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=7; refFlag[7]=0;  end 
14'h1244: begin refPos[0]=2; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=0; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=2; refFlag[6]=0; refPos[7]=3; refFlag[7]=0;  end 
14'h1245: begin refPos[0]=6; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=0; refFlag[6]=1; refPos[7]=99; refFlag[7]=2;  end 
14'h1246: begin refPos[0]=10; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=4; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h1247: begin refPos[0]=14; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=8; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h1250: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=23; refFlag[7]=0;  end 
14'h1251: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=19; refFlag[7]=0;  end 
14'h1252: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=15; refFlag[7]=0;  end 
14'h1253: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=11; refFlag[7]=0;  end 
14'h1254: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=7; refFlag[7]=0;  end 
14'h1255: begin refPos[0]=2; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=0; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=2; refFlag[6]=0; refPos[7]=3; refFlag[7]=0;  end 
14'h1256: begin refPos[0]=6; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=0; refFlag[6]=1; refPos[7]=99; refFlag[7]=2;  end 
14'h1257: begin refPos[0]=10; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=4; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h1260: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=26; refFlag[6]=0; refPos[7]=27; refFlag[7]=0;  end 
14'h1261: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=23; refFlag[7]=0;  end 
14'h1262: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=19; refFlag[7]=0;  end 
14'h1263: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=15; refFlag[7]=0;  end 
14'h1264: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=11; refFlag[7]=0;  end 
14'h1265: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=7; refFlag[7]=0;  end 
14'h1266: begin refPos[0]=2; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=0; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=2; refFlag[6]=0; refPos[7]=3; refFlag[7]=0;  end 
14'h1267: begin refPos[0]=6; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=0; refFlag[6]=1; refPos[7]=99; refFlag[7]=2;  end 
14'h1270: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=30; refFlag[6]=0; refPos[7]=31; refFlag[7]=0;  end 
14'h1271: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=26; refFlag[6]=0; refPos[7]=27; refFlag[7]=0;  end 
14'h1272: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=23; refFlag[7]=0;  end 
14'h1273: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=19; refFlag[7]=0;  end 
14'h1274: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=15; refFlag[7]=0;  end 
14'h1275: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=11; refFlag[7]=0;  end 
14'h1276: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=7; refFlag[7]=0;  end 
14'h1277: begin refPos[0]=2; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=0; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=2; refFlag[6]=0; refPos[7]=3; refFlag[7]=0;  end 
14'h1300: begin refPos[0]=3; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=0; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=2; refFlag[6]=0; refPos[7]=3; refFlag[7]=0;  end 
14'h1301: begin refPos[0]=6; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=0; refFlag[5]=1; refPos[6]=99; refFlag[6]=2; refPos[7]=0; refFlag[7]=0;  end 
14'h1302: begin refPos[0]=10; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=3; refFlag[6]=1; refPos[7]=1; refFlag[7]=1;  end 
14'h1303: begin refPos[0]=14; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=5; refFlag[7]=1;  end 
14'h1304: begin refPos[0]=19; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=15; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=10; refFlag[7]=1;  end 
14'h1305: begin refPos[0]=22; refFlag[0]=1; refPos[1]=21; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=15; refFlag[6]=1; refPos[7]=14; refFlag[7]=1;  end 
14'h1306: begin refPos[0]=26; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=21; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=19; refFlag[6]=1; refPos[7]=17; refFlag[7]=1;  end 
14'h1307: begin refPos[0]=30; refFlag[0]=1; refPos[1]=29; refFlag[1]=1; refPos[2]=27; refFlag[2]=1; refPos[3]=26; refFlag[3]=1; refPos[4]=25; refFlag[4]=1; refPos[5]=24; refFlag[5]=1; refPos[6]=22; refFlag[6]=1; refPos[7]=21; refFlag[7]=1;  end 
14'h1310: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=7; refFlag[7]=0;  end 
14'h1311: begin refPos[0]=1; refFlag[0]=1; refPos[1]=0; refFlag[1]=1; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=2; refFlag[5]=0; refPos[6]=3; refFlag[6]=0; refPos[7]=4; refFlag[7]=0;  end 
14'h1312: begin refPos[0]=5; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=0; refFlag[4]=1; refPos[5]=99; refFlag[5]=2; refPos[6]=0; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h1313: begin refPos[0]=9; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=3; refFlag[5]=1; refPos[6]=1; refFlag[6]=1; refPos[7]=0; refFlag[7]=1;  end 
14'h1314: begin refPos[0]=14; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=5; refFlag[7]=1;  end 
14'h1315: begin refPos[0]=17; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=15; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=9; refFlag[7]=1;  end 
14'h1316: begin refPos[0]=21; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=15; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=13; refFlag[7]=1;  end 
14'h1317: begin refPos[0]=25; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=16; refFlag[7]=1;  end 
14'h1320: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=11; refFlag[7]=0;  end 
14'h1321: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=7; refFlag[6]=0; refPos[7]=8; refFlag[7]=0;  end 
14'h1322: begin refPos[0]=0; refFlag[0]=1; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=2; refFlag[4]=0; refPos[5]=3; refFlag[5]=0; refPos[6]=4; refFlag[6]=0; refPos[7]=5; refFlag[7]=0;  end 
14'h1323: begin refPos[0]=4; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=0; refFlag[3]=1; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=2; refFlag[7]=0;  end 
14'h1324: begin refPos[0]=9; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=3; refFlag[5]=1; refPos[6]=1; refFlag[6]=1; refPos[7]=0; refFlag[7]=1;  end 
14'h1325: begin refPos[0]=13; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=5; refFlag[6]=1; refPos[7]=4; refFlag[7]=1;  end 
14'h1326: begin refPos[0]=16; refFlag[0]=1; refPos[1]=15; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=9; refFlag[6]=1; refPos[7]=8; refFlag[7]=1;  end 
14'h1327: begin refPos[0]=20; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=15; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=13; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h1330: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=15; refFlag[7]=0;  end 
14'h1331: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=12; refFlag[7]=0;  end 
14'h1332: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=8; refFlag[6]=0; refPos[7]=9; refFlag[7]=0;  end 
14'h1333: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=5; refFlag[6]=0; refPos[7]=6; refFlag[7]=0;  end 
14'h1334: begin refPos[0]=4; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=0; refFlag[3]=1; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=2; refFlag[7]=0;  end 
14'h1335: begin refPos[0]=8; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=0; refFlag[6]=1; refPos[7]=99; refFlag[7]=2;  end 
14'h1336: begin refPos[0]=11; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=4; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h1337: begin refPos[0]=15; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=8; refFlag[6]=1; refPos[7]=6; refFlag[7]=1;  end 
14'h1340: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=19; refFlag[7]=0;  end 
14'h1341: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=15; refFlag[6]=0; refPos[7]=16; refFlag[7]=0;  end 
14'h1342: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=12; refFlag[6]=0; refPos[7]=13; refFlag[7]=0;  end 
14'h1343: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=9; refFlag[6]=0; refPos[7]=10; refFlag[7]=0;  end 
14'h1344: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=5; refFlag[6]=0; refPos[7]=6; refFlag[7]=0;  end 
14'h1345: begin refPos[0]=3; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=0; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=2; refFlag[6]=0; refPos[7]=3; refFlag[7]=0;  end 
14'h1346: begin refPos[0]=6; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=0; refFlag[5]=1; refPos[6]=99; refFlag[6]=2; refPos[7]=0; refFlag[7]=0;  end 
14'h1347: begin refPos[0]=10; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=3; refFlag[6]=1; refPos[7]=1; refFlag[7]=1;  end 
14'h1350: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=23; refFlag[7]=0;  end 
14'h1351: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=20; refFlag[7]=0;  end 
14'h1352: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=16; refFlag[6]=0; refPos[7]=17; refFlag[7]=0;  end 
14'h1353: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=13; refFlag[6]=0; refPos[7]=14; refFlag[7]=0;  end 
14'h1354: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=9; refFlag[6]=0; refPos[7]=10; refFlag[7]=0;  end 
14'h1355: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=7; refFlag[7]=0;  end 
14'h1356: begin refPos[0]=1; refFlag[0]=1; refPos[1]=0; refFlag[1]=1; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=2; refFlag[5]=0; refPos[6]=3; refFlag[6]=0; refPos[7]=4; refFlag[7]=0;  end 
14'h1357: begin refPos[0]=5; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=0; refFlag[4]=1; refPos[5]=99; refFlag[5]=2; refPos[6]=0; refFlag[6]=0; refPos[7]=1; refFlag[7]=0;  end 
14'h1360: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=26; refFlag[6]=0; refPos[7]=27; refFlag[7]=0;  end 
14'h1361: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=24; refFlag[7]=0;  end 
14'h1362: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=20; refFlag[6]=0; refPos[7]=21; refFlag[7]=0;  end 
14'h1363: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=18; refFlag[7]=0;  end 
14'h1364: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=13; refFlag[6]=0; refPos[7]=14; refFlag[7]=0;  end 
14'h1365: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=11; refFlag[7]=0;  end 
14'h1366: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=7; refFlag[6]=0; refPos[7]=8; refFlag[7]=0;  end 
14'h1367: begin refPos[0]=0; refFlag[0]=1; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=2; refFlag[4]=0; refPos[5]=3; refFlag[5]=0; refPos[6]=4; refFlag[6]=0; refPos[7]=5; refFlag[7]=0;  end 
14'h1370: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=30; refFlag[6]=0; refPos[7]=31; refFlag[7]=0;  end 
14'h1371: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=28; refFlag[7]=0;  end 
14'h1372: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=24; refFlag[6]=0; refPos[7]=25; refFlag[7]=0;  end 
14'h1373: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=21; refFlag[6]=0; refPos[7]=22; refFlag[7]=0;  end 
14'h1374: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=18; refFlag[7]=0;  end 
14'h1375: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=15; refFlag[7]=0;  end 
14'h1376: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=12; refFlag[7]=0;  end 
14'h1377: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=8; refFlag[6]=0; refPos[7]=9; refFlag[7]=0;  end 
14'h1400: begin refPos[0]=2; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=2; refFlag[5]=0; refPos[6]=3; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1401: begin refPos[0]=7; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=99; refFlag[5]=2; refPos[6]=0; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1402: begin refPos[0]=10; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=2; refFlag[5]=1; refPos[6]=1; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1403: begin refPos[0]=14; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=5; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1404: begin refPos[0]=19; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=11; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1405: begin refPos[0]=22; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=19; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=13; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1406: begin refPos[0]=26; refFlag[0]=1; refPos[1]=25; refFlag[1]=1; refPos[2]=23; refFlag[2]=1; refPos[3]=22; refFlag[3]=1; refPos[4]=20; refFlag[4]=1; refPos[5]=19; refFlag[5]=1; refPos[6]=17; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1407: begin refPos[0]=29; refFlag[0]=1; refPos[1]=28; refFlag[1]=1; refPos[2]=26; refFlag[2]=1; refPos[3]=25; refFlag[3]=1; refPos[4]=23; refFlag[4]=1; refPos[5]=22; refFlag[5]=1; refPos[6]=20; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1410: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=7; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1411: begin refPos[0]=1; refFlag[0]=1; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=2; refFlag[4]=0; refPos[5]=3; refFlag[5]=0; refPos[6]=4; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1412: begin refPos[0]=4; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=2; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1413: begin refPos[0]=8; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=99; refFlag[6]=2; refPos[7]=1; refFlag[7]=-1;  end 
14'h1414: begin refPos[0]=13; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=4; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1415: begin refPos[0]=16; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=7; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1416: begin refPos[0]=20; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1417: begin refPos[0]=23; refFlag[0]=1; refPos[1]=22; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=17; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1420: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1421: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=8; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1422: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1423: begin refPos[0]=2; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=2; refFlag[5]=0; refPos[6]=3; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1424: begin refPos[0]=7; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=2; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=99; refFlag[5]=2; refPos[6]=0; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1425: begin refPos[0]=10; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=2; refFlag[5]=1; refPos[6]=1; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1426: begin refPos[0]=14; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=8; refFlag[4]=1; refPos[5]=7; refFlag[5]=1; refPos[6]=5; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1427: begin refPos[0]=17; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=8; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1430: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=15; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1431: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=12; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1432: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1433: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=7; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1434: begin refPos[0]=1; refFlag[0]=1; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=2; refFlag[4]=0; refPos[5]=3; refFlag[5]=0; refPos[6]=4; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1435: begin refPos[0]=4; refFlag[0]=1; refPos[1]=2; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=2; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1436: begin refPos[0]=8; refFlag[0]=1; refPos[1]=7; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=2; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=99; refFlag[6]=2; refPos[7]=1; refFlag[7]=-1;  end 
14'h1437: begin refPos[0]=11; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=8; refFlag[2]=1; refPos[3]=7; refFlag[3]=1; refPos[4]=5; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1440: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1441: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=16; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1442: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1443: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1444: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=8; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1445: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1446: begin refPos[0]=2; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=2; refFlag[5]=0; refPos[6]=3; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1447: begin refPos[0]=5; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=2; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1450: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1451: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=20; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1452: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1453: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=15; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1454: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=12; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1455: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1456: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=7; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1457: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=5; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1460: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1461: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=24; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1462: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1463: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1464: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=16; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1465: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1466: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1467: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=9; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1470: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=31; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1471: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=27; refFlag[5]=0; refPos[6]=28; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1472: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=26; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1473: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1474: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=20; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1475: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1476: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=15; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1477: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=13; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1500: begin refPos[0]=3; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=2; refFlag[5]=0; refPos[6]=3; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1501: begin refPos[0]=7; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1502: begin refPos[0]=10; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=99; refFlag[6]=2; refPos[7]=1; refFlag[7]=-1;  end 
14'h1503: begin refPos[0]=14; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=3; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1504: begin refPos[0]=18; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=7; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1505: begin refPos[0]=22; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1506: begin refPos[0]=25; refFlag[0]=1; refPos[1]=23; refFlag[1]=1; refPos[2]=22; refFlag[2]=1; refPos[3]=20; refFlag[3]=1; refPos[4]=18; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1507: begin refPos[0]=29; refFlag[0]=1; refPos[1]=27; refFlag[1]=1; refPos[2]=25; refFlag[2]=1; refPos[3]=23; refFlag[3]=1; refPos[4]=22; refFlag[4]=1; refPos[5]=20; refFlag[5]=1; refPos[6]=18; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1510: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=7; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1511: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=5; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1512: begin refPos[0]=3; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=2; refFlag[5]=0; refPos[6]=3; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1513: begin refPos[0]=7; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1514: begin refPos[0]=10; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=99; refFlag[6]=2; refPos[7]=1; refFlag[7]=-1;  end 
14'h1515: begin refPos[0]=14; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=3; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1516: begin refPos[0]=18; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=12; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=8; refFlag[5]=1; refPos[6]=7; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1517: begin refPos[0]=22; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=18; refFlag[2]=1; refPos[3]=16; refFlag[3]=1; refPos[4]=14; refFlag[4]=1; refPos[5]=12; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1520: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1521: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=9; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1522: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=7; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1523: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=5; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1524: begin refPos[0]=3; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=2; refFlag[5]=0; refPos[6]=3; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1525: begin refPos[0]=7; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1526: begin refPos[0]=10; refFlag[0]=1; refPos[1]=8; refFlag[1]=1; refPos[2]=7; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=99; refFlag[6]=2; refPos[7]=1; refFlag[7]=-1;  end 
14'h1527: begin refPos[0]=14; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=8; refFlag[3]=1; refPos[4]=7; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=3; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1530: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=15; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1531: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=13; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1532: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1533: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=9; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1534: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=7; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1535: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=5; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1536: begin refPos[0]=3; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=2; refFlag[5]=0; refPos[6]=3; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1537: begin refPos[0]=7; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1540: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1541: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1542: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=15; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1543: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=13; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1544: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1545: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=9; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1546: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=7; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1547: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=5; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1550: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1551: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=21; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1552: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1553: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1554: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=15; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1555: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=13; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1556: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1557: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=9; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1560: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1561: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=25; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1562: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1563: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=21; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1564: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1565: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1566: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=15; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1567: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=13; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1570: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=31; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1571: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=29; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1572: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1573: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=25; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1574: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1575: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=21; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1576: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1577: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1600: begin refPos[0]=1; refFlag[0]=1; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=2; refFlag[4]=0; refPos[5]=3; refFlag[5]=0; refPos[6]=4; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1601: begin refPos[0]=6; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=2; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1602: begin refPos[0]=9; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1603: begin refPos[0]=14; refFlag[0]=1; refPos[1]=11; refFlag[1]=1; refPos[2]=9; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=4; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=99; refFlag[6]=2; refPos[7]=1; refFlag[7]=-1;  end 
14'h1604: begin refPos[0]=19; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=4; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1605: begin refPos[0]=21; refFlag[0]=1; refPos[1]=19; refFlag[1]=1; refPos[2]=16; refFlag[2]=1; refPos[3]=14; refFlag[3]=1; refPos[4]=11; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1606: begin refPos[0]=26; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=21; refFlag[2]=1; refPos[3]=19; refFlag[3]=1; refPos[4]=16; refFlag[4]=1; refPos[5]=14; refFlag[5]=1; refPos[6]=11; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1607: begin refPos[0]=29; refFlag[0]=1; refPos[1]=26; refFlag[1]=1; refPos[2]=24; refFlag[2]=1; refPos[3]=21; refFlag[3]=1; refPos[4]=19; refFlag[4]=1; refPos[5]=16; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1610: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=8; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1611: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1612: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=5; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1613: begin refPos[0]=4; refFlag[0]=1; refPos[1]=1; refFlag[1]=1; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=2; refFlag[5]=0; refPos[6]=3; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1614: begin refPos[0]=9; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1615: begin refPos[0]=11; refFlag[0]=1; refPos[1]=9; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=4; refFlag[3]=1; refPos[4]=1; refFlag[4]=1; refPos[5]=99; refFlag[5]=2; refPos[6]=0; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1616: begin refPos[0]=16; refFlag[0]=1; refPos[1]=14; refFlag[1]=1; refPos[2]=11; refFlag[2]=1; refPos[3]=9; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=4; refFlag[5]=1; refPos[6]=1; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1617: begin refPos[0]=19; refFlag[0]=1; refPos[1]=16; refFlag[1]=1; refPos[2]=14; refFlag[2]=1; refPos[3]=11; refFlag[3]=1; refPos[4]=9; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=4; refFlag[6]=1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1620: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=12; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1621: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1622: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=9; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1623: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=7; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1624: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=5; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1625: begin refPos[0]=1; refFlag[0]=1; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=2; refFlag[4]=0; refPos[5]=3; refFlag[5]=0; refPos[6]=4; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1626: begin refPos[0]=6; refFlag[0]=1; refPos[1]=4; refFlag[1]=1; refPos[2]=1; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=2; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1627: begin refPos[0]=9; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=4; refFlag[2]=1; refPos[3]=1; refFlag[3]=1; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=0; refPos[6]=1; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1630: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=16; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1631: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1632: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=13; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1633: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1634: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=9; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1635: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=8; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1636: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1637: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=5; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1640: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=20; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1641: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1642: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1643: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=15; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1644: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=13; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1645: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=12; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1646: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1647: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=9; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1650: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=24; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1651: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1652: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=21; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1653: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1654: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1655: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=16; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1656: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1657: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=13; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1660: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=27; refFlag[5]=0; refPos[6]=28; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1661: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=26; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1662: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=25; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1663: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1664: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=21; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1665: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=20; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1666: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1667: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1670: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=31; refFlag[5]=0; refPos[6]=32; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1671: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=30; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1672: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=29; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1673: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1674: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=25; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1675: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=24; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1676: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1677: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=21; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1700: begin refPos[0]=3; refFlag[0]=1; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=2; refFlag[4]=0; refPos[5]=3; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1701: begin refPos[0]=6; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=2; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1702: begin refPos[0]=10; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1703: begin refPos[0]=13; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1704: begin refPos[0]=17; refFlag[0]=1; refPos[1]=13; refFlag[1]=1; refPos[2]=10; refFlag[2]=1; refPos[3]=6; refFlag[3]=1; refPos[4]=3; refFlag[4]=1; refPos[5]=99; refFlag[5]=2; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1705: begin refPos[0]=20; refFlag[0]=1; refPos[1]=17; refFlag[1]=1; refPos[2]=13; refFlag[2]=1; refPos[3]=10; refFlag[3]=1; refPos[4]=6; refFlag[4]=1; refPos[5]=3; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1706: begin refPos[0]=24; refFlag[0]=1; refPos[1]=20; refFlag[1]=1; refPos[2]=17; refFlag[2]=1; refPos[3]=13; refFlag[3]=1; refPos[4]=10; refFlag[4]=1; refPos[5]=6; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1707: begin refPos[0]=27; refFlag[0]=1; refPos[1]=24; refFlag[1]=1; refPos[2]=20; refFlag[2]=1; refPos[3]=17; refFlag[3]=1; refPos[4]=13; refFlag[4]=1; refPos[5]=10; refFlag[5]=1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1710: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1711: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1712: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1713: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1714: begin refPos[0]=3; refFlag[0]=1; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=2; refFlag[4]=0; refPos[5]=3; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1715: begin refPos[0]=6; refFlag[0]=1; refPos[1]=3; refFlag[1]=1; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=2; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1716: begin refPos[0]=10; refFlag[0]=1; refPos[1]=6; refFlag[1]=1; refPos[2]=3; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1717: begin refPos[0]=13; refFlag[0]=1; refPos[1]=10; refFlag[1]=1; refPos[2]=6; refFlag[2]=1; refPos[3]=3; refFlag[3]=1; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1720: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1721: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1722: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1723: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1724: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1725: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1726: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1727: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1730: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1731: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1732: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1733: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1734: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1735: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1736: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1737: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1740: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1741: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1742: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1743: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1744: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1745: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1746: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1747: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1750: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1751: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1752: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1753: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1754: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1755: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1756: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1757: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1760: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=27; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1761: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1762: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1763: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1764: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1765: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1766: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1767: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1770: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=31; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1771: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1772: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1773: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1774: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=27; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1775: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1776: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1777: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1800: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1801: begin refPos[0]=5; refFlag[0]=1; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=2; refFlag[4]=0; refPos[5]=3; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1802: begin refPos[0]=5; refFlag[0]=1; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=2; refFlag[4]=0; refPos[5]=3; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1803: begin refPos[0]=12; refFlag[0]=1; refPos[1]=5; refFlag[1]=1; refPos[2]=99; refFlag[2]=2; refPos[3]=0; refFlag[3]=0; refPos[4]=1; refFlag[4]=0; refPos[5]=2; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1804: begin refPos[0]=18; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1805: begin refPos[0]=18; refFlag[0]=1; refPos[1]=12; refFlag[1]=1; refPos[2]=5; refFlag[2]=1; refPos[3]=99; refFlag[3]=2; refPos[4]=0; refFlag[4]=0; refPos[5]=1; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1806: begin refPos[0]=25; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1807: begin refPos[0]=25; refFlag[0]=1; refPos[1]=18; refFlag[1]=1; refPos[2]=12; refFlag[2]=1; refPos[3]=5; refFlag[3]=1; refPos[4]=99; refFlag[4]=2; refPos[5]=0; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1810: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1811: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1812: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1813: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1814: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1815: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1816: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1817: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=4; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1820: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1821: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1822: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1823: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1824: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1825: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1826: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1827: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1830: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1831: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1832: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1833: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1834: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1835: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1836: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1837: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1840: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1841: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1842: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1843: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1844: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1845: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1846: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1847: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1850: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1851: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1852: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1853: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1854: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1855: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1856: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1857: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1860: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1861: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=27; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1862: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=27; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1863: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1864: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1865: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1866: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1867: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1870: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=32; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1871: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=31; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1872: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=31; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1873: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1874: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1875: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1876: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1877: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1900: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1901: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1902: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1903: begin refPos[0]=99; refFlag[0]=2; refPos[1]=0; refFlag[1]=0; refPos[2]=1; refFlag[2]=0; refPos[3]=2; refFlag[3]=0; refPos[4]=3; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1904: begin refPos[0]=15; refFlag[0]=1; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=2; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1905: begin refPos[0]=15; refFlag[0]=1; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=2; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1906: begin refPos[0]=15; refFlag[0]=1; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=2; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1907: begin refPos[0]=15; refFlag[0]=1; refPos[1]=99; refFlag[1]=2; refPos[2]=0; refFlag[2]=0; refPos[3]=1; refFlag[3]=0; refPos[4]=2; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1910: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1911: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1912: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1913: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1914: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1915: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1916: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1917: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1920: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1921: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1922: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1923: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1924: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1925: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1926: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1927: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1930: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1931: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1932: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1933: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1934: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1935: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1936: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1937: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1940: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1941: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1942: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1943: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1944: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1945: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1946: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1947: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1950: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1951: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1952: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1953: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1954: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1955: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1956: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1957: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1960: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1961: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1962: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1963: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1964: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1965: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1966: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1967: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1970: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1971: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1972: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1973: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1974: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1975: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1976: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1977: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a00: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=0; refFlag[4]=1; refPos[5]=1; refFlag[5]=1; refPos[6]=2; refFlag[6]=1; refPos[7]=3; refFlag[7]=1;  end 
14'h1a01: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=1; refPos[5]=5; refFlag[5]=1; refPos[6]=6; refFlag[6]=1; refPos[7]=7; refFlag[7]=1;  end 
14'h1a02: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=8; refFlag[4]=1; refPos[5]=9; refFlag[5]=1; refPos[6]=10; refFlag[6]=1; refPos[7]=11; refFlag[7]=1;  end 
14'h1a03: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=12; refFlag[4]=1; refPos[5]=13; refFlag[5]=1; refPos[6]=14; refFlag[6]=1; refPos[7]=15; refFlag[7]=1;  end 
14'h1a04: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a05: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a06: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a07: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a10: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a11: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a12: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a13: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a14: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a15: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a16: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a17: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a20: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a21: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a22: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a23: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a24: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a25: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a26: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a27: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a30: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a31: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a32: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a33: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a34: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a35: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a36: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a37: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a40: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a41: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a42: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a43: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a44: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a45: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a46: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a47: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a50: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a51: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a52: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a53: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a54: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a55: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a56: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a57: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a60: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a61: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a62: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a63: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a64: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a65: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a66: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a67: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a70: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a71: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a72: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a73: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a74: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a75: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a76: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1a77: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=1; refFlag[4]=-1; refPos[5]=1; refFlag[5]=-1; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b00: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b01: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b02: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b03: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b04: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b05: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b06: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b07: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b10: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b11: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b12: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b13: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b14: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b15: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b16: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b17: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b20: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b21: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b22: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b23: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b24: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b25: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b26: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b27: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b30: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b31: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b32: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b33: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b34: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b35: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b36: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b37: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b40: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b41: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b42: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b43: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b44: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b45: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b46: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b47: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b50: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b51: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b52: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b53: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b54: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b55: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b56: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b57: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b60: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b61: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b62: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b63: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b64: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b65: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b66: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b67: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b70: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b71: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b72: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b73: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b74: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b75: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b76: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1b77: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c00: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c01: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c02: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c03: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c04: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c05: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c06: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c07: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c10: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c11: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c12: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c13: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c14: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c15: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c16: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c17: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c20: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c21: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c22: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c23: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c24: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c25: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c26: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c27: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c30: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c31: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c32: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c33: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c34: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c35: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c36: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c37: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c40: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c41: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c42: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c43: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c44: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c45: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c46: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c47: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c50: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c51: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c52: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c53: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=27; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c54: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=27; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c55: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c56: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c57: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c60: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c61: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c62: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c63: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=31; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c64: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=31; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c65: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=32; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c66: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=32; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c67: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c70: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c71: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c72: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c73: begin refPos[0]=30; refFlag[0]=0; refPos[1]=31; refFlag[1]=0; refPos[2]=32; refFlag[2]=0; refPos[3]=33; refFlag[3]=0; refPos[4]=34; refFlag[4]=0; refPos[5]=35; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c74: begin refPos[0]=30; refFlag[0]=0; refPos[1]=31; refFlag[1]=0; refPos[2]=32; refFlag[2]=0; refPos[3]=33; refFlag[3]=0; refPos[4]=34; refFlag[4]=0; refPos[5]=35; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c75: begin refPos[0]=31; refFlag[0]=0; refPos[1]=32; refFlag[1]=0; refPos[2]=33; refFlag[2]=0; refPos[3]=34; refFlag[3]=0; refPos[4]=35; refFlag[4]=0; refPos[5]=36; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c76: begin refPos[0]=31; refFlag[0]=0; refPos[1]=32; refFlag[1]=0; refPos[2]=33; refFlag[2]=0; refPos[3]=34; refFlag[3]=0; refPos[4]=35; refFlag[4]=0; refPos[5]=36; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1c77: begin refPos[0]=32; refFlag[0]=0; refPos[1]=33; refFlag[1]=0; refPos[2]=34; refFlag[2]=0; refPos[3]=35; refFlag[3]=0; refPos[4]=36; refFlag[4]=0; refPos[5]=37; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d00: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d01: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d02: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d03: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d04: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d05: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d06: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d07: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d10: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d11: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d12: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d13: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d14: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d15: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d16: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d17: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d20: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d21: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d22: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d23: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d24: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d25: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d26: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d27: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d30: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d31: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d32: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d33: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d34: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d35: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d36: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d37: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d40: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d41: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d42: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d43: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d44: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d45: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d46: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d47: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d50: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d51: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d52: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=27; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d53: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d54: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d55: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d56: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=32; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d57: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d60: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d61: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d62: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=31; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d63: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=32; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d64: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d65: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d66: begin refPos[0]=31; refFlag[0]=0; refPos[1]=32; refFlag[1]=0; refPos[2]=33; refFlag[2]=0; refPos[3]=34; refFlag[3]=0; refPos[4]=35; refFlag[4]=0; refPos[5]=36; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d67: begin refPos[0]=32; refFlag[0]=0; refPos[1]=33; refFlag[1]=0; refPos[2]=34; refFlag[2]=0; refPos[3]=35; refFlag[3]=0; refPos[4]=36; refFlag[4]=0; refPos[5]=37; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d70: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d71: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d72: begin refPos[0]=30; refFlag[0]=0; refPos[1]=31; refFlag[1]=0; refPos[2]=32; refFlag[2]=0; refPos[3]=33; refFlag[3]=0; refPos[4]=34; refFlag[4]=0; refPos[5]=35; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d73: begin refPos[0]=31; refFlag[0]=0; refPos[1]=32; refFlag[1]=0; refPos[2]=33; refFlag[2]=0; refPos[3]=34; refFlag[3]=0; refPos[4]=35; refFlag[4]=0; refPos[5]=36; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d74: begin refPos[0]=32; refFlag[0]=0; refPos[1]=33; refFlag[1]=0; refPos[2]=34; refFlag[2]=0; refPos[3]=35; refFlag[3]=0; refPos[4]=36; refFlag[4]=0; refPos[5]=37; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d75: begin refPos[0]=33; refFlag[0]=0; refPos[1]=34; refFlag[1]=0; refPos[2]=35; refFlag[2]=0; refPos[3]=36; refFlag[3]=0; refPos[4]=37; refFlag[4]=0; refPos[5]=38; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d76: begin refPos[0]=35; refFlag[0]=0; refPos[1]=36; refFlag[1]=0; refPos[2]=37; refFlag[2]=0; refPos[3]=38; refFlag[3]=0; refPos[4]=39; refFlag[4]=0; refPos[5]=40; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1d77: begin refPos[0]=36; refFlag[0]=0; refPos[1]=37; refFlag[1]=0; refPos[2]=38; refFlag[2]=0; refPos[3]=39; refFlag[3]=0; refPos[4]=40; refFlag[4]=0; refPos[5]=41; refFlag[5]=0; refPos[6]=1; refFlag[6]=-1; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e00: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e01: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=8; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e02: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=9; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e03: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e04: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=12; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e05: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e06: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=16; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e07: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e10: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e11: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=12; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e12: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=13; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e13: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=15; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e14: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=16; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e15: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e16: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=20; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e17: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=21; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e20: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e21: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=16; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e22: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e23: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e24: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=20; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e25: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e26: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=24; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e27: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=25; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e30: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e31: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=20; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e32: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=21; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e33: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e34: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=24; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e35: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=26; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e36: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=27; refFlag[5]=0; refPos[6]=28; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e37: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=29; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e40: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e41: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=24; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e42: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=25; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e43: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e44: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=27; refFlag[5]=0; refPos[6]=28; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e45: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=30; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e46: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=31; refFlag[5]=0; refPos[6]=32; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e47: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=32; refFlag[5]=0; refPos[6]=33; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e50: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=26; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e51: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=27; refFlag[5]=0; refPos[6]=28; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e52: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=29; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e53: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=31; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e54: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=31; refFlag[5]=0; refPos[6]=32; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e55: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=34; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e56: begin refPos[0]=30; refFlag[0]=0; refPos[1]=31; refFlag[1]=0; refPos[2]=32; refFlag[2]=0; refPos[3]=33; refFlag[3]=0; refPos[4]=34; refFlag[4]=0; refPos[5]=35; refFlag[5]=0; refPos[6]=36; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e57: begin refPos[0]=31; refFlag[0]=0; refPos[1]=32; refFlag[1]=0; refPos[2]=33; refFlag[2]=0; refPos[3]=34; refFlag[3]=0; refPos[4]=35; refFlag[4]=0; refPos[5]=36; refFlag[5]=0; refPos[6]=37; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e60: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=30; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e61: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=31; refFlag[5]=0; refPos[6]=32; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e62: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=32; refFlag[5]=0; refPos[6]=33; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e63: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=35; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e64: begin refPos[0]=30; refFlag[0]=0; refPos[1]=31; refFlag[1]=0; refPos[2]=32; refFlag[2]=0; refPos[3]=33; refFlag[3]=0; refPos[4]=34; refFlag[4]=0; refPos[5]=35; refFlag[5]=0; refPos[6]=36; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e65: begin refPos[0]=32; refFlag[0]=0; refPos[1]=33; refFlag[1]=0; refPos[2]=34; refFlag[2]=0; refPos[3]=35; refFlag[3]=0; refPos[4]=36; refFlag[4]=0; refPos[5]=37; refFlag[5]=0; refPos[6]=38; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e66: begin refPos[0]=34; refFlag[0]=0; refPos[1]=35; refFlag[1]=0; refPos[2]=36; refFlag[2]=0; refPos[3]=37; refFlag[3]=0; refPos[4]=38; refFlag[4]=0; refPos[5]=39; refFlag[5]=0; refPos[6]=40; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e67: begin refPos[0]=35; refFlag[0]=0; refPos[1]=36; refFlag[1]=0; refPos[2]=37; refFlag[2]=0; refPos[3]=38; refFlag[3]=0; refPos[4]=39; refFlag[4]=0; refPos[5]=40; refFlag[5]=0; refPos[6]=41; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e70: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=34; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e71: begin refPos[0]=30; refFlag[0]=0; refPos[1]=31; refFlag[1]=0; refPos[2]=32; refFlag[2]=0; refPos[3]=33; refFlag[3]=0; refPos[4]=34; refFlag[4]=0; refPos[5]=35; refFlag[5]=0; refPos[6]=36; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e72: begin refPos[0]=31; refFlag[0]=0; refPos[1]=32; refFlag[1]=0; refPos[2]=33; refFlag[2]=0; refPos[3]=34; refFlag[3]=0; refPos[4]=35; refFlag[4]=0; refPos[5]=36; refFlag[5]=0; refPos[6]=37; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e73: begin refPos[0]=33; refFlag[0]=0; refPos[1]=34; refFlag[1]=0; refPos[2]=35; refFlag[2]=0; refPos[3]=36; refFlag[3]=0; refPos[4]=37; refFlag[4]=0; refPos[5]=38; refFlag[5]=0; refPos[6]=39; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e74: begin refPos[0]=34; refFlag[0]=0; refPos[1]=35; refFlag[1]=0; refPos[2]=36; refFlag[2]=0; refPos[3]=37; refFlag[3]=0; refPos[4]=38; refFlag[4]=0; refPos[5]=39; refFlag[5]=0; refPos[6]=40; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e75: begin refPos[0]=36; refFlag[0]=0; refPos[1]=37; refFlag[1]=0; refPos[2]=38; refFlag[2]=0; refPos[3]=39; refFlag[3]=0; refPos[4]=40; refFlag[4]=0; refPos[5]=41; refFlag[5]=0; refPos[6]=42; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e76: begin refPos[0]=38; refFlag[0]=0; refPos[1]=39; refFlag[1]=0; refPos[2]=40; refFlag[2]=0; refPos[3]=41; refFlag[3]=0; refPos[4]=42; refFlag[4]=0; refPos[5]=43; refFlag[5]=0; refPos[6]=44; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1e77: begin refPos[0]=39; refFlag[0]=0; refPos[1]=40; refFlag[1]=0; refPos[2]=41; refFlag[2]=0; refPos[3]=42; refFlag[3]=0; refPos[4]=43; refFlag[4]=0; refPos[5]=44; refFlag[5]=0; refPos[6]=45; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f00: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f01: begin refPos[0]=2; refFlag[0]=0; refPos[1]=3; refFlag[1]=0; refPos[2]=4; refFlag[2]=0; refPos[3]=5; refFlag[3]=0; refPos[4]=6; refFlag[4]=0; refPos[5]=7; refFlag[5]=0; refPos[6]=8; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f02: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f03: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=12; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f04: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=15; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f05: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f06: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f07: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=21; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f10: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f11: begin refPos[0]=6; refFlag[0]=0; refPos[1]=7; refFlag[1]=0; refPos[2]=8; refFlag[2]=0; refPos[3]=9; refFlag[3]=0; refPos[4]=10; refFlag[4]=0; refPos[5]=11; refFlag[5]=0; refPos[6]=12; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f12: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f13: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=16; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f14: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f15: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=21; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f16: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f17: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=25; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f20: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f21: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=16; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f22: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f23: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=20; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f24: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f25: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=25; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f26: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f27: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=29; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f30: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f31: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=20; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f32: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f33: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=24; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f34: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f35: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=29; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f36: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=31; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f37: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=32; refFlag[5]=0; refPos[6]=33; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f40: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f41: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=24; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f42: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=26; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f43: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=27; refFlag[5]=0; refPos[6]=28; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f44: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=31; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f45: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=32; refFlag[5]=0; refPos[6]=33; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f46: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=35; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f47: begin refPos[0]=31; refFlag[0]=0; refPos[1]=32; refFlag[1]=0; refPos[2]=33; refFlag[2]=0; refPos[3]=34; refFlag[3]=0; refPos[4]=35; refFlag[4]=0; refPos[5]=36; refFlag[5]=0; refPos[6]=37; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f50: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=26; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f51: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=27; refFlag[5]=0; refPos[6]=28; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f52: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=30; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f53: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=31; refFlag[5]=0; refPos[6]=32; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f54: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=35; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f55: begin refPos[0]=31; refFlag[0]=0; refPos[1]=32; refFlag[1]=0; refPos[2]=33; refFlag[2]=0; refPos[3]=34; refFlag[3]=0; refPos[4]=35; refFlag[4]=0; refPos[5]=36; refFlag[5]=0; refPos[6]=37; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f56: begin refPos[0]=33; refFlag[0]=0; refPos[1]=34; refFlag[1]=0; refPos[2]=35; refFlag[2]=0; refPos[3]=36; refFlag[3]=0; refPos[4]=37; refFlag[4]=0; refPos[5]=38; refFlag[5]=0; refPos[6]=39; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f57: begin refPos[0]=35; refFlag[0]=0; refPos[1]=36; refFlag[1]=0; refPos[2]=37; refFlag[2]=0; refPos[3]=38; refFlag[3]=0; refPos[4]=39; refFlag[4]=0; refPos[5]=40; refFlag[5]=0; refPos[6]=41; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f60: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=30; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f61: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=31; refFlag[5]=0; refPos[6]=32; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f62: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=34; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f63: begin refPos[0]=30; refFlag[0]=0; refPos[1]=31; refFlag[1]=0; refPos[2]=32; refFlag[2]=0; refPos[3]=33; refFlag[3]=0; refPos[4]=34; refFlag[4]=0; refPos[5]=35; refFlag[5]=0; refPos[6]=36; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f64: begin refPos[0]=33; refFlag[0]=0; refPos[1]=34; refFlag[1]=0; refPos[2]=35; refFlag[2]=0; refPos[3]=36; refFlag[3]=0; refPos[4]=37; refFlag[4]=0; refPos[5]=38; refFlag[5]=0; refPos[6]=39; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f65: begin refPos[0]=35; refFlag[0]=0; refPos[1]=36; refFlag[1]=0; refPos[2]=37; refFlag[2]=0; refPos[3]=38; refFlag[3]=0; refPos[4]=39; refFlag[4]=0; refPos[5]=40; refFlag[5]=0; refPos[6]=41; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f66: begin refPos[0]=37; refFlag[0]=0; refPos[1]=38; refFlag[1]=0; refPos[2]=39; refFlag[2]=0; refPos[3]=40; refFlag[3]=0; refPos[4]=41; refFlag[4]=0; refPos[5]=42; refFlag[5]=0; refPos[6]=43; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f67: begin refPos[0]=39; refFlag[0]=0; refPos[1]=40; refFlag[1]=0; refPos[2]=41; refFlag[2]=0; refPos[3]=42; refFlag[3]=0; refPos[4]=43; refFlag[4]=0; refPos[5]=44; refFlag[5]=0; refPos[6]=45; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f70: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=34; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f71: begin refPos[0]=30; refFlag[0]=0; refPos[1]=31; refFlag[1]=0; refPos[2]=32; refFlag[2]=0; refPos[3]=33; refFlag[3]=0; refPos[4]=34; refFlag[4]=0; refPos[5]=35; refFlag[5]=0; refPos[6]=36; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f72: begin refPos[0]=32; refFlag[0]=0; refPos[1]=33; refFlag[1]=0; refPos[2]=34; refFlag[2]=0; refPos[3]=35; refFlag[3]=0; refPos[4]=36; refFlag[4]=0; refPos[5]=37; refFlag[5]=0; refPos[6]=38; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f73: begin refPos[0]=34; refFlag[0]=0; refPos[1]=35; refFlag[1]=0; refPos[2]=36; refFlag[2]=0; refPos[3]=37; refFlag[3]=0; refPos[4]=38; refFlag[4]=0; refPos[5]=39; refFlag[5]=0; refPos[6]=40; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f74: begin refPos[0]=37; refFlag[0]=0; refPos[1]=38; refFlag[1]=0; refPos[2]=39; refFlag[2]=0; refPos[3]=40; refFlag[3]=0; refPos[4]=41; refFlag[4]=0; refPos[5]=42; refFlag[5]=0; refPos[6]=43; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f75: begin refPos[0]=39; refFlag[0]=0; refPos[1]=40; refFlag[1]=0; refPos[2]=41; refFlag[2]=0; refPos[3]=42; refFlag[3]=0; refPos[4]=43; refFlag[4]=0; refPos[5]=44; refFlag[5]=0; refPos[6]=45; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f76: begin refPos[0]=41; refFlag[0]=0; refPos[1]=42; refFlag[1]=0; refPos[2]=43; refFlag[2]=0; refPos[3]=44; refFlag[3]=0; refPos[4]=45; refFlag[4]=0; refPos[5]=46; refFlag[5]=0; refPos[6]=47; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h1f77: begin refPos[0]=43; refFlag[0]=0; refPos[1]=44; refFlag[1]=0; refPos[2]=45; refFlag[2]=0; refPos[3]=46; refFlag[3]=0; refPos[4]=47; refFlag[4]=0; refPos[5]=48; refFlag[5]=0; refPos[6]=49; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2000: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2001: begin refPos[0]=3; refFlag[0]=0; refPos[1]=4; refFlag[1]=0; refPos[2]=5; refFlag[2]=0; refPos[3]=6; refFlag[3]=0; refPos[4]=7; refFlag[4]=0; refPos[5]=8; refFlag[5]=0; refPos[6]=9; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2002: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2003: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2004: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2005: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2006: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2007: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=25; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2010: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2011: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=13; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2012: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=15; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2013: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2014: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=21; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2015: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2016: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=26; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2017: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=29; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2020: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2021: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2022: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2023: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2024: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=25; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2025: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2026: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=30; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2027: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=32; refFlag[5]=0; refPos[6]=33; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2030: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2031: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=21; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2032: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2033: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=26; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2034: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=29; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2035: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=31; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2036: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=34; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2037: begin refPos[0]=31; refFlag[0]=0; refPos[1]=32; refFlag[1]=0; refPos[2]=33; refFlag[2]=0; refPos[3]=34; refFlag[3]=0; refPos[4]=35; refFlag[4]=0; refPos[5]=36; refFlag[5]=0; refPos[6]=37; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2040: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2041: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=25; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2042: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2043: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=30; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2044: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=32; refFlag[5]=0; refPos[6]=33; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2045: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=35; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2046: begin refPos[0]=32; refFlag[0]=0; refPos[1]=33; refFlag[1]=0; refPos[2]=34; refFlag[2]=0; refPos[3]=35; refFlag[3]=0; refPos[4]=36; refFlag[4]=0; refPos[5]=37; refFlag[5]=0; refPos[6]=38; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2047: begin refPos[0]=35; refFlag[0]=0; refPos[1]=36; refFlag[1]=0; refPos[2]=37; refFlag[2]=0; refPos[3]=38; refFlag[3]=0; refPos[4]=39; refFlag[4]=0; refPos[5]=40; refFlag[5]=0; refPos[6]=41; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2050: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=26; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2051: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=29; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2052: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=31; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2053: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=34; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2054: begin refPos[0]=31; refFlag[0]=0; refPos[1]=32; refFlag[1]=0; refPos[2]=33; refFlag[2]=0; refPos[3]=34; refFlag[3]=0; refPos[4]=35; refFlag[4]=0; refPos[5]=36; refFlag[5]=0; refPos[6]=37; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2055: begin refPos[0]=33; refFlag[0]=0; refPos[1]=34; refFlag[1]=0; refPos[2]=35; refFlag[2]=0; refPos[3]=36; refFlag[3]=0; refPos[4]=37; refFlag[4]=0; refPos[5]=38; refFlag[5]=0; refPos[6]=39; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2056: begin refPos[0]=36; refFlag[0]=0; refPos[1]=37; refFlag[1]=0; refPos[2]=38; refFlag[2]=0; refPos[3]=39; refFlag[3]=0; refPos[4]=40; refFlag[4]=0; refPos[5]=41; refFlag[5]=0; refPos[6]=42; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2057: begin refPos[0]=39; refFlag[0]=0; refPos[1]=40; refFlag[1]=0; refPos[2]=41; refFlag[2]=0; refPos[3]=42; refFlag[3]=0; refPos[4]=43; refFlag[4]=0; refPos[5]=44; refFlag[5]=0; refPos[6]=45; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2060: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=30; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2061: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=32; refFlag[5]=0; refPos[6]=33; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2062: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=35; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2063: begin refPos[0]=32; refFlag[0]=0; refPos[1]=33; refFlag[1]=0; refPos[2]=34; refFlag[2]=0; refPos[3]=35; refFlag[3]=0; refPos[4]=36; refFlag[4]=0; refPos[5]=37; refFlag[5]=0; refPos[6]=38; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2064: begin refPos[0]=35; refFlag[0]=0; refPos[1]=36; refFlag[1]=0; refPos[2]=37; refFlag[2]=0; refPos[3]=38; refFlag[3]=0; refPos[4]=39; refFlag[4]=0; refPos[5]=40; refFlag[5]=0; refPos[6]=41; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2065: begin refPos[0]=37; refFlag[0]=0; refPos[1]=38; refFlag[1]=0; refPos[2]=39; refFlag[2]=0; refPos[3]=40; refFlag[3]=0; refPos[4]=41; refFlag[4]=0; refPos[5]=42; refFlag[5]=0; refPos[6]=43; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2066: begin refPos[0]=40; refFlag[0]=0; refPos[1]=41; refFlag[1]=0; refPos[2]=42; refFlag[2]=0; refPos[3]=43; refFlag[3]=0; refPos[4]=44; refFlag[4]=0; refPos[5]=45; refFlag[5]=0; refPos[6]=46; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2067: begin refPos[0]=43; refFlag[0]=0; refPos[1]=44; refFlag[1]=0; refPos[2]=45; refFlag[2]=0; refPos[3]=46; refFlag[3]=0; refPos[4]=47; refFlag[4]=0; refPos[5]=48; refFlag[5]=0; refPos[6]=49; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2070: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=34; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2071: begin refPos[0]=31; refFlag[0]=0; refPos[1]=32; refFlag[1]=0; refPos[2]=33; refFlag[2]=0; refPos[3]=34; refFlag[3]=0; refPos[4]=35; refFlag[4]=0; refPos[5]=36; refFlag[5]=0; refPos[6]=37; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2072: begin refPos[0]=33; refFlag[0]=0; refPos[1]=34; refFlag[1]=0; refPos[2]=35; refFlag[2]=0; refPos[3]=36; refFlag[3]=0; refPos[4]=37; refFlag[4]=0; refPos[5]=38; refFlag[5]=0; refPos[6]=39; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2073: begin refPos[0]=36; refFlag[0]=0; refPos[1]=37; refFlag[1]=0; refPos[2]=38; refFlag[2]=0; refPos[3]=39; refFlag[3]=0; refPos[4]=40; refFlag[4]=0; refPos[5]=41; refFlag[5]=0; refPos[6]=42; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2074: begin refPos[0]=39; refFlag[0]=0; refPos[1]=40; refFlag[1]=0; refPos[2]=41; refFlag[2]=0; refPos[3]=42; refFlag[3]=0; refPos[4]=43; refFlag[4]=0; refPos[5]=44; refFlag[5]=0; refPos[6]=45; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2075: begin refPos[0]=41; refFlag[0]=0; refPos[1]=42; refFlag[1]=0; refPos[2]=43; refFlag[2]=0; refPos[3]=44; refFlag[3]=0; refPos[4]=45; refFlag[4]=0; refPos[5]=46; refFlag[5]=0; refPos[6]=47; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2076: begin refPos[0]=44; refFlag[0]=0; refPos[1]=45; refFlag[1]=0; refPos[2]=46; refFlag[2]=0; refPos[3]=47; refFlag[3]=0; refPos[4]=48; refFlag[4]=0; refPos[5]=49; refFlag[5]=0; refPos[6]=50; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2077: begin refPos[0]=47; refFlag[0]=0; refPos[1]=48; refFlag[1]=0; refPos[2]=49; refFlag[2]=0; refPos[3]=50; refFlag[3]=0; refPos[4]=51; refFlag[4]=0; refPos[5]=52; refFlag[5]=0; refPos[6]=53; refFlag[6]=0; refPos[7]=1; refFlag[7]=-1;  end 
14'h2100: begin refPos[0]=0; refFlag[0]=0; refPos[1]=1; refFlag[1]=0; refPos[2]=2; refFlag[2]=0; refPos[3]=3; refFlag[3]=0; refPos[4]=4; refFlag[4]=0; refPos[5]=5; refFlag[5]=0; refPos[6]=6; refFlag[6]=0; refPos[7]=7; refFlag[7]=0;  end 
14'h2101: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=11; refFlag[7]=0;  end 
14'h2102: begin refPos[0]=7; refFlag[0]=0; refPos[1]=8; refFlag[1]=0; refPos[2]=9; refFlag[2]=0; refPos[3]=10; refFlag[3]=0; refPos[4]=11; refFlag[4]=0; refPos[5]=12; refFlag[5]=0; refPos[6]=13; refFlag[6]=0; refPos[7]=14; refFlag[7]=0;  end 
14'h2103: begin refPos[0]=10; refFlag[0]=0; refPos[1]=11; refFlag[1]=0; refPos[2]=12; refFlag[2]=0; refPos[3]=13; refFlag[3]=0; refPos[4]=14; refFlag[4]=0; refPos[5]=15; refFlag[5]=0; refPos[6]=16; refFlag[6]=0; refPos[7]=17; refFlag[7]=0;  end 
14'h2104: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=20; refFlag[7]=0;  end 
14'h2105: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=24; refFlag[7]=0;  end 
14'h2106: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=26; refFlag[6]=0; refPos[7]=27; refFlag[7]=0;  end 
14'h2107: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=29; refFlag[6]=0; refPos[7]=30; refFlag[7]=0;  end 
14'h2110: begin refPos[0]=4; refFlag[0]=0; refPos[1]=5; refFlag[1]=0; refPos[2]=6; refFlag[2]=0; refPos[3]=7; refFlag[3]=0; refPos[4]=8; refFlag[4]=0; refPos[5]=9; refFlag[5]=0; refPos[6]=10; refFlag[6]=0; refPos[7]=11; refFlag[7]=0;  end 
14'h2111: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=15; refFlag[7]=0;  end 
14'h2112: begin refPos[0]=11; refFlag[0]=0; refPos[1]=12; refFlag[1]=0; refPos[2]=13; refFlag[2]=0; refPos[3]=14; refFlag[3]=0; refPos[4]=15; refFlag[4]=0; refPos[5]=16; refFlag[5]=0; refPos[6]=17; refFlag[6]=0; refPos[7]=18; refFlag[7]=0;  end 
14'h2113: begin refPos[0]=14; refFlag[0]=0; refPos[1]=15; refFlag[1]=0; refPos[2]=16; refFlag[2]=0; refPos[3]=17; refFlag[3]=0; refPos[4]=18; refFlag[4]=0; refPos[5]=19; refFlag[5]=0; refPos[6]=20; refFlag[6]=0; refPos[7]=21; refFlag[7]=0;  end 
14'h2114: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=24; refFlag[7]=0;  end 
14'h2115: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=28; refFlag[7]=0;  end 
14'h2116: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=30; refFlag[6]=0; refPos[7]=31; refFlag[7]=0;  end 
14'h2117: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=32; refFlag[5]=0; refPos[6]=33; refFlag[6]=0; refPos[7]=34; refFlag[7]=0;  end 
14'h2120: begin refPos[0]=8; refFlag[0]=0; refPos[1]=9; refFlag[1]=0; refPos[2]=10; refFlag[2]=0; refPos[3]=11; refFlag[3]=0; refPos[4]=12; refFlag[4]=0; refPos[5]=13; refFlag[5]=0; refPos[6]=14; refFlag[6]=0; refPos[7]=15; refFlag[7]=0;  end 
14'h2121: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=19; refFlag[7]=0;  end 
14'h2122: begin refPos[0]=15; refFlag[0]=0; refPos[1]=16; refFlag[1]=0; refPos[2]=17; refFlag[2]=0; refPos[3]=18; refFlag[3]=0; refPos[4]=19; refFlag[4]=0; refPos[5]=20; refFlag[5]=0; refPos[6]=21; refFlag[6]=0; refPos[7]=22; refFlag[7]=0;  end 
14'h2123: begin refPos[0]=18; refFlag[0]=0; refPos[1]=19; refFlag[1]=0; refPos[2]=20; refFlag[2]=0; refPos[3]=21; refFlag[3]=0; refPos[4]=22; refFlag[4]=0; refPos[5]=23; refFlag[5]=0; refPos[6]=24; refFlag[6]=0; refPos[7]=25; refFlag[7]=0;  end 
14'h2124: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=28; refFlag[7]=0;  end 
14'h2125: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=31; refFlag[6]=0; refPos[7]=32; refFlag[7]=0;  end 
14'h2126: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=34; refFlag[6]=0; refPos[7]=35; refFlag[7]=0;  end 
14'h2127: begin refPos[0]=31; refFlag[0]=0; refPos[1]=32; refFlag[1]=0; refPos[2]=33; refFlag[2]=0; refPos[3]=34; refFlag[3]=0; refPos[4]=35; refFlag[4]=0; refPos[5]=36; refFlag[5]=0; refPos[6]=37; refFlag[6]=0; refPos[7]=38; refFlag[7]=0;  end 
14'h2130: begin refPos[0]=12; refFlag[0]=0; refPos[1]=13; refFlag[1]=0; refPos[2]=14; refFlag[2]=0; refPos[3]=15; refFlag[3]=0; refPos[4]=16; refFlag[4]=0; refPos[5]=17; refFlag[5]=0; refPos[6]=18; refFlag[6]=0; refPos[7]=19; refFlag[7]=0;  end 
14'h2131: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=23; refFlag[7]=0;  end 
14'h2132: begin refPos[0]=19; refFlag[0]=0; refPos[1]=20; refFlag[1]=0; refPos[2]=21; refFlag[2]=0; refPos[3]=22; refFlag[3]=0; refPos[4]=23; refFlag[4]=0; refPos[5]=24; refFlag[5]=0; refPos[6]=25; refFlag[6]=0; refPos[7]=26; refFlag[7]=0;  end 
14'h2133: begin refPos[0]=22; refFlag[0]=0; refPos[1]=23; refFlag[1]=0; refPos[2]=24; refFlag[2]=0; refPos[3]=25; refFlag[3]=0; refPos[4]=26; refFlag[4]=0; refPos[5]=27; refFlag[5]=0; refPos[6]=28; refFlag[6]=0; refPos[7]=29; refFlag[7]=0;  end 
14'h2134: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=31; refFlag[6]=0; refPos[7]=32; refFlag[7]=0;  end 
14'h2135: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=35; refFlag[6]=0; refPos[7]=36; refFlag[7]=0;  end 
14'h2136: begin refPos[0]=32; refFlag[0]=0; refPos[1]=33; refFlag[1]=0; refPos[2]=34; refFlag[2]=0; refPos[3]=35; refFlag[3]=0; refPos[4]=36; refFlag[4]=0; refPos[5]=37; refFlag[5]=0; refPos[6]=38; refFlag[6]=0; refPos[7]=39; refFlag[7]=0;  end 
14'h2137: begin refPos[0]=35; refFlag[0]=0; refPos[1]=36; refFlag[1]=0; refPos[2]=37; refFlag[2]=0; refPos[3]=38; refFlag[3]=0; refPos[4]=39; refFlag[4]=0; refPos[5]=40; refFlag[5]=0; refPos[6]=41; refFlag[6]=0; refPos[7]=42; refFlag[7]=0;  end 
14'h2140: begin refPos[0]=16; refFlag[0]=0; refPos[1]=17; refFlag[1]=0; refPos[2]=18; refFlag[2]=0; refPos[3]=19; refFlag[3]=0; refPos[4]=20; refFlag[4]=0; refPos[5]=21; refFlag[5]=0; refPos[6]=22; refFlag[6]=0; refPos[7]=23; refFlag[7]=0;  end 
14'h2141: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=26; refFlag[6]=0; refPos[7]=27; refFlag[7]=0;  end 
14'h2142: begin refPos[0]=23; refFlag[0]=0; refPos[1]=24; refFlag[1]=0; refPos[2]=25; refFlag[2]=0; refPos[3]=26; refFlag[3]=0; refPos[4]=27; refFlag[4]=0; refPos[5]=28; refFlag[5]=0; refPos[6]=29; refFlag[6]=0; refPos[7]=30; refFlag[7]=0;  end 
14'h2143: begin refPos[0]=26; refFlag[0]=0; refPos[1]=27; refFlag[1]=0; refPos[2]=28; refFlag[2]=0; refPos[3]=29; refFlag[3]=0; refPos[4]=30; refFlag[4]=0; refPos[5]=31; refFlag[5]=0; refPos[6]=32; refFlag[6]=0; refPos[7]=33; refFlag[7]=0;  end 
14'h2144: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=35; refFlag[6]=0; refPos[7]=36; refFlag[7]=0;  end 
14'h2145: begin refPos[0]=33; refFlag[0]=0; refPos[1]=34; refFlag[1]=0; refPos[2]=35; refFlag[2]=0; refPos[3]=36; refFlag[3]=0; refPos[4]=37; refFlag[4]=0; refPos[5]=38; refFlag[5]=0; refPos[6]=39; refFlag[6]=0; refPos[7]=40; refFlag[7]=0;  end 
14'h2146: begin refPos[0]=36; refFlag[0]=0; refPos[1]=37; refFlag[1]=0; refPos[2]=38; refFlag[2]=0; refPos[3]=39; refFlag[3]=0; refPos[4]=40; refFlag[4]=0; refPos[5]=41; refFlag[5]=0; refPos[6]=42; refFlag[6]=0; refPos[7]=43; refFlag[7]=0;  end 
14'h2147: begin refPos[0]=39; refFlag[0]=0; refPos[1]=40; refFlag[1]=0; refPos[2]=41; refFlag[2]=0; refPos[3]=42; refFlag[3]=0; refPos[4]=43; refFlag[4]=0; refPos[5]=44; refFlag[5]=0; refPos[6]=45; refFlag[6]=0; refPos[7]=46; refFlag[7]=0;  end 
14'h2150: begin refPos[0]=20; refFlag[0]=0; refPos[1]=21; refFlag[1]=0; refPos[2]=22; refFlag[2]=0; refPos[3]=23; refFlag[3]=0; refPos[4]=24; refFlag[4]=0; refPos[5]=25; refFlag[5]=0; refPos[6]=26; refFlag[6]=0; refPos[7]=27; refFlag[7]=0;  end 
14'h2151: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=30; refFlag[6]=0; refPos[7]=31; refFlag[7]=0;  end 
14'h2152: begin refPos[0]=27; refFlag[0]=0; refPos[1]=28; refFlag[1]=0; refPos[2]=29; refFlag[2]=0; refPos[3]=30; refFlag[3]=0; refPos[4]=31; refFlag[4]=0; refPos[5]=32; refFlag[5]=0; refPos[6]=33; refFlag[6]=0; refPos[7]=34; refFlag[7]=0;  end 
14'h2153: begin refPos[0]=30; refFlag[0]=0; refPos[1]=31; refFlag[1]=0; refPos[2]=32; refFlag[2]=0; refPos[3]=33; refFlag[3]=0; refPos[4]=34; refFlag[4]=0; refPos[5]=35; refFlag[5]=0; refPos[6]=36; refFlag[6]=0; refPos[7]=37; refFlag[7]=0;  end 
14'h2154: begin refPos[0]=33; refFlag[0]=0; refPos[1]=34; refFlag[1]=0; refPos[2]=35; refFlag[2]=0; refPos[3]=36; refFlag[3]=0; refPos[4]=37; refFlag[4]=0; refPos[5]=38; refFlag[5]=0; refPos[6]=39; refFlag[6]=0; refPos[7]=40; refFlag[7]=0;  end 
14'h2155: begin refPos[0]=37; refFlag[0]=0; refPos[1]=38; refFlag[1]=0; refPos[2]=39; refFlag[2]=0; refPos[3]=40; refFlag[3]=0; refPos[4]=41; refFlag[4]=0; refPos[5]=42; refFlag[5]=0; refPos[6]=43; refFlag[6]=0; refPos[7]=44; refFlag[7]=0;  end 
14'h2156: begin refPos[0]=40; refFlag[0]=0; refPos[1]=41; refFlag[1]=0; refPos[2]=42; refFlag[2]=0; refPos[3]=43; refFlag[3]=0; refPos[4]=44; refFlag[4]=0; refPos[5]=45; refFlag[5]=0; refPos[6]=46; refFlag[6]=0; refPos[7]=47; refFlag[7]=0;  end 
14'h2157: begin refPos[0]=43; refFlag[0]=0; refPos[1]=44; refFlag[1]=0; refPos[2]=45; refFlag[2]=0; refPos[3]=46; refFlag[3]=0; refPos[4]=47; refFlag[4]=0; refPos[5]=48; refFlag[5]=0; refPos[6]=49; refFlag[6]=0; refPos[7]=50; refFlag[7]=0;  end 
14'h2160: begin refPos[0]=24; refFlag[0]=0; refPos[1]=25; refFlag[1]=0; refPos[2]=26; refFlag[2]=0; refPos[3]=27; refFlag[3]=0; refPos[4]=28; refFlag[4]=0; refPos[5]=29; refFlag[5]=0; refPos[6]=30; refFlag[6]=0; refPos[7]=31; refFlag[7]=0;  end 
14'h2161: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=34; refFlag[6]=0; refPos[7]=35; refFlag[7]=0;  end 
14'h2162: begin refPos[0]=31; refFlag[0]=0; refPos[1]=32; refFlag[1]=0; refPos[2]=33; refFlag[2]=0; refPos[3]=34; refFlag[3]=0; refPos[4]=35; refFlag[4]=0; refPos[5]=36; refFlag[5]=0; refPos[6]=37; refFlag[6]=0; refPos[7]=38; refFlag[7]=0;  end 
14'h2163: begin refPos[0]=34; refFlag[0]=0; refPos[1]=35; refFlag[1]=0; refPos[2]=36; refFlag[2]=0; refPos[3]=37; refFlag[3]=0; refPos[4]=38; refFlag[4]=0; refPos[5]=39; refFlag[5]=0; refPos[6]=40; refFlag[6]=0; refPos[7]=41; refFlag[7]=0;  end 
14'h2164: begin refPos[0]=37; refFlag[0]=0; refPos[1]=38; refFlag[1]=0; refPos[2]=39; refFlag[2]=0; refPos[3]=40; refFlag[3]=0; refPos[4]=41; refFlag[4]=0; refPos[5]=42; refFlag[5]=0; refPos[6]=43; refFlag[6]=0; refPos[7]=44; refFlag[7]=0;  end 
14'h2165: begin refPos[0]=41; refFlag[0]=0; refPos[1]=42; refFlag[1]=0; refPos[2]=43; refFlag[2]=0; refPos[3]=44; refFlag[3]=0; refPos[4]=45; refFlag[4]=0; refPos[5]=46; refFlag[5]=0; refPos[6]=47; refFlag[6]=0; refPos[7]=48; refFlag[7]=0;  end 
14'h2166: begin refPos[0]=44; refFlag[0]=0; refPos[1]=45; refFlag[1]=0; refPos[2]=46; refFlag[2]=0; refPos[3]=47; refFlag[3]=0; refPos[4]=48; refFlag[4]=0; refPos[5]=49; refFlag[5]=0; refPos[6]=50; refFlag[6]=0; refPos[7]=51; refFlag[7]=0;  end 
14'h2167: begin refPos[0]=47; refFlag[0]=0; refPos[1]=48; refFlag[1]=0; refPos[2]=49; refFlag[2]=0; refPos[3]=50; refFlag[3]=0; refPos[4]=51; refFlag[4]=0; refPos[5]=52; refFlag[5]=0; refPos[6]=53; refFlag[6]=0; refPos[7]=54; refFlag[7]=0;  end 
14'h2170: begin refPos[0]=28; refFlag[0]=0; refPos[1]=29; refFlag[1]=0; refPos[2]=30; refFlag[2]=0; refPos[3]=31; refFlag[3]=0; refPos[4]=32; refFlag[4]=0; refPos[5]=33; refFlag[5]=0; refPos[6]=34; refFlag[6]=0; refPos[7]=35; refFlag[7]=0;  end 
14'h2171: begin refPos[0]=32; refFlag[0]=0; refPos[1]=33; refFlag[1]=0; refPos[2]=34; refFlag[2]=0; refPos[3]=35; refFlag[3]=0; refPos[4]=36; refFlag[4]=0; refPos[5]=37; refFlag[5]=0; refPos[6]=38; refFlag[6]=0; refPos[7]=39; refFlag[7]=0;  end 
14'h2172: begin refPos[0]=35; refFlag[0]=0; refPos[1]=36; refFlag[1]=0; refPos[2]=37; refFlag[2]=0; refPos[3]=38; refFlag[3]=0; refPos[4]=39; refFlag[4]=0; refPos[5]=40; refFlag[5]=0; refPos[6]=41; refFlag[6]=0; refPos[7]=42; refFlag[7]=0;  end 
14'h2173: begin refPos[0]=38; refFlag[0]=0; refPos[1]=39; refFlag[1]=0; refPos[2]=40; refFlag[2]=0; refPos[3]=41; refFlag[3]=0; refPos[4]=42; refFlag[4]=0; refPos[5]=43; refFlag[5]=0; refPos[6]=44; refFlag[6]=0; refPos[7]=45; refFlag[7]=0;  end 
14'h2174: begin refPos[0]=41; refFlag[0]=0; refPos[1]=42; refFlag[1]=0; refPos[2]=43; refFlag[2]=0; refPos[3]=44; refFlag[3]=0; refPos[4]=45; refFlag[4]=0; refPos[5]=46; refFlag[5]=0; refPos[6]=47; refFlag[6]=0; refPos[7]=48; refFlag[7]=0;  end 
14'h2175: begin refPos[0]=45; refFlag[0]=0; refPos[1]=46; refFlag[1]=0; refPos[2]=47; refFlag[2]=0; refPos[3]=48; refFlag[3]=0; refPos[4]=49; refFlag[4]=0; refPos[5]=50; refFlag[5]=0; refPos[6]=51; refFlag[6]=0; refPos[7]=52; refFlag[7]=0;  end 
14'h2176: begin refPos[0]=48; refFlag[0]=0; refPos[1]=49; refFlag[1]=0; refPos[2]=50; refFlag[2]=0; refPos[3]=51; refFlag[3]=0; refPos[4]=52; refFlag[4]=0; refPos[5]=53; refFlag[5]=0; refPos[6]=54; refFlag[6]=0; refPos[7]=55; refFlag[7]=0;  end 
14'h2177: begin refPos[0]=51; refFlag[0]=0; refPos[1]=52; refFlag[1]=0; refPos[2]=53; refFlag[2]=0; refPos[3]=54; refFlag[3]=0; refPos[4]=55; refFlag[4]=0; refPos[5]=56; refFlag[5]=0; refPos[6]=57; refFlag[6]=0; refPos[7]=58; refFlag[7]=0;  end 
14'h2200: begin refPos[0]=1; refFlag[0]=0; refPos[1]=2; refFlag[1]=0; refPos[2]=3; refFlag[2]=0; refPos[3]=4; refFlag[3]=0; refPos[4]=5; refFlag[4]=0; refPos[5]=6; refFlag[5]=0; refPos[6]=7; refFlag[6]=0; if(tuSize!=2) refPos[7]=8; else refPos[7]=7; refFlag[7]=0;  end 
14'h2201: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=12; refFlag[7]=0;  end 
14'h2202: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=15; refFlag[6]=0; refPos[7]=16; refFlag[7]=0;  end 
14'h2203: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=20; refFlag[7]=0;  end 
14'h2204: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=24; refFlag[7]=0;  end 
14'h2205: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=28; refFlag[7]=0;  end 
14'h2206: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=31; refFlag[6]=0; refPos[7]=32; refFlag[7]=0;  end 
14'h2207: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=35; refFlag[6]=0; refPos[7]=36; refFlag[7]=0;  end 
14'h2210: begin refPos[0]=5; refFlag[0]=0; refPos[1]=6; refFlag[1]=0; refPos[2]=7; refFlag[2]=0; refPos[3]=8; refFlag[3]=0; refPos[4]=9; refFlag[4]=0; refPos[5]=10; refFlag[5]=0; refPos[6]=11; refFlag[6]=0; refPos[7]=12; refFlag[7]=0;  end 
14'h2211: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=15; refFlag[6]=0; if(tuSize!=3)refPos[7]=16; else refPos[7]=15; refFlag[7]=0;  end 
14'h2212: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=20; refFlag[7]=0;  end 
14'h2213: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=24; refFlag[7]=0;  end 
14'h2214: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=28; refFlag[7]=0;  end 
14'h2215: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=31; refFlag[6]=0; refPos[7]=32; refFlag[7]=0;  end 
14'h2216: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=35; refFlag[6]=0; refPos[7]=36; refFlag[7]=0;  end 
14'h2217: begin refPos[0]=33; refFlag[0]=0; refPos[1]=34; refFlag[1]=0; refPos[2]=35; refFlag[2]=0; refPos[3]=36; refFlag[3]=0; refPos[4]=37; refFlag[4]=0; refPos[5]=38; refFlag[5]=0; refPos[6]=39; refFlag[6]=0; refPos[7]=40; refFlag[7]=0;  end 
14'h2220: begin refPos[0]=9; refFlag[0]=0; refPos[1]=10; refFlag[1]=0; refPos[2]=11; refFlag[2]=0; refPos[3]=12; refFlag[3]=0; refPos[4]=13; refFlag[4]=0; refPos[5]=14; refFlag[5]=0; refPos[6]=15; refFlag[6]=0; refPos[7]=16; refFlag[7]=0;  end 
14'h2221: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=20; refFlag[7]=0;  end 
14'h2222: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=24; refFlag[7]=0;  end 
14'h2223: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=28; refFlag[7]=0;  end 
14'h2224: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=31; refFlag[6]=0; refPos[7]=32; refFlag[7]=0;  end 
14'h2225: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=35; refFlag[6]=0; refPos[7]=36; refFlag[7]=0;  end 
14'h2226: begin refPos[0]=33; refFlag[0]=0; refPos[1]=34; refFlag[1]=0; refPos[2]=35; refFlag[2]=0; refPos[3]=36; refFlag[3]=0; refPos[4]=37; refFlag[4]=0; refPos[5]=38; refFlag[5]=0; refPos[6]=39; refFlag[6]=0; refPos[7]=40; refFlag[7]=0;  end 
14'h2227: begin refPos[0]=37; refFlag[0]=0; refPos[1]=38; refFlag[1]=0; refPos[2]=39; refFlag[2]=0; refPos[3]=40; refFlag[3]=0; refPos[4]=41; refFlag[4]=0; refPos[5]=42; refFlag[5]=0; refPos[6]=43; refFlag[6]=0; refPos[7]=44; refFlag[7]=0;  end 
14'h2230: begin refPos[0]=13; refFlag[0]=0; refPos[1]=14; refFlag[1]=0; refPos[2]=15; refFlag[2]=0; refPos[3]=16; refFlag[3]=0; refPos[4]=17; refFlag[4]=0; refPos[5]=18; refFlag[5]=0; refPos[6]=19; refFlag[6]=0; refPos[7]=20; refFlag[7]=0;  end 
14'h2231: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=24; refFlag[7]=0;  end 
14'h2232: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=28; refFlag[7]=0;  end 
14'h2233: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=31; refFlag[6]=0; if(tuSize!=4) refPos[7]=32; else refPos[7]=31; refFlag[7]=0;  end 
14'h2234: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=35; refFlag[6]=0; refPos[7]=36; refFlag[7]=0;  end 
14'h2235: begin refPos[0]=33; refFlag[0]=0; refPos[1]=34; refFlag[1]=0; refPos[2]=35; refFlag[2]=0; refPos[3]=36; refFlag[3]=0; refPos[4]=37; refFlag[4]=0; refPos[5]=38; refFlag[5]=0; refPos[6]=39; refFlag[6]=0; refPos[7]=40; refFlag[7]=0;  end 
14'h2236: begin refPos[0]=37; refFlag[0]=0; refPos[1]=38; refFlag[1]=0; refPos[2]=39; refFlag[2]=0; refPos[3]=40; refFlag[3]=0; refPos[4]=41; refFlag[4]=0; refPos[5]=42; refFlag[5]=0; refPos[6]=43; refFlag[6]=0; refPos[7]=44; refFlag[7]=0;  end 
14'h2237: begin refPos[0]=41; refFlag[0]=0; refPos[1]=42; refFlag[1]=0; refPos[2]=43; refFlag[2]=0; refPos[3]=44; refFlag[3]=0; refPos[4]=45; refFlag[4]=0; refPos[5]=46; refFlag[5]=0; refPos[6]=47; refFlag[6]=0; refPos[7]=48; refFlag[7]=0;  end 
14'h2240: begin refPos[0]=17; refFlag[0]=0; refPos[1]=18; refFlag[1]=0; refPos[2]=19; refFlag[2]=0; refPos[3]=20; refFlag[3]=0; refPos[4]=21; refFlag[4]=0; refPos[5]=22; refFlag[5]=0; refPos[6]=23; refFlag[6]=0; refPos[7]=24; refFlag[7]=0;  end 
14'h2241: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=28; refFlag[7]=0;  end 
14'h2242: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=31; refFlag[6]=0; refPos[7]=32; refFlag[7]=0;  end 
14'h2243: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=35; refFlag[6]=0; refPos[7]=36; refFlag[7]=0;  end 
14'h2244: begin refPos[0]=33; refFlag[0]=0; refPos[1]=34; refFlag[1]=0; refPos[2]=35; refFlag[2]=0; refPos[3]=36; refFlag[3]=0; refPos[4]=37; refFlag[4]=0; refPos[5]=38; refFlag[5]=0; refPos[6]=39; refFlag[6]=0; refPos[7]=40; refFlag[7]=0;  end 
14'h2245: begin refPos[0]=37; refFlag[0]=0; refPos[1]=38; refFlag[1]=0; refPos[2]=39; refFlag[2]=0; refPos[3]=40; refFlag[3]=0; refPos[4]=41; refFlag[4]=0; refPos[5]=42; refFlag[5]=0; refPos[6]=43; refFlag[6]=0; refPos[7]=44; refFlag[7]=0;  end 
14'h2246: begin refPos[0]=41; refFlag[0]=0; refPos[1]=42; refFlag[1]=0; refPos[2]=43; refFlag[2]=0; refPos[3]=44; refFlag[3]=0; refPos[4]=45; refFlag[4]=0; refPos[5]=46; refFlag[5]=0; refPos[6]=47; refFlag[6]=0; refPos[7]=48; refFlag[7]=0;  end 
14'h2247: begin refPos[0]=45; refFlag[0]=0; refPos[1]=46; refFlag[1]=0; refPos[2]=47; refFlag[2]=0; refPos[3]=48; refFlag[3]=0; refPos[4]=49; refFlag[4]=0; refPos[5]=50; refFlag[5]=0; refPos[6]=51; refFlag[6]=0; refPos[7]=52; refFlag[7]=0;  end 
14'h2250: begin refPos[0]=21; refFlag[0]=0; refPos[1]=22; refFlag[1]=0; refPos[2]=23; refFlag[2]=0; refPos[3]=24; refFlag[3]=0; refPos[4]=25; refFlag[4]=0; refPos[5]=26; refFlag[5]=0; refPos[6]=27; refFlag[6]=0; refPos[7]=28; refFlag[7]=0;  end 
14'h2251: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=31; refFlag[6]=0; refPos[7]=32; refFlag[7]=0;  end 
14'h2252: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=35; refFlag[6]=0; refPos[7]=36; refFlag[7]=0;  end 
14'h2253: begin refPos[0]=33; refFlag[0]=0; refPos[1]=34; refFlag[1]=0; refPos[2]=35; refFlag[2]=0; refPos[3]=36; refFlag[3]=0; refPos[4]=37; refFlag[4]=0; refPos[5]=38; refFlag[5]=0; refPos[6]=39; refFlag[6]=0; refPos[7]=40; refFlag[7]=0;  end 
14'h2254: begin refPos[0]=37; refFlag[0]=0; refPos[1]=38; refFlag[1]=0; refPos[2]=39; refFlag[2]=0; refPos[3]=40; refFlag[3]=0; refPos[4]=41; refFlag[4]=0; refPos[5]=42; refFlag[5]=0; refPos[6]=43; refFlag[6]=0; refPos[7]=44; refFlag[7]=0;  end 
14'h2255: begin refPos[0]=41; refFlag[0]=0; refPos[1]=42; refFlag[1]=0; refPos[2]=43; refFlag[2]=0; refPos[3]=44; refFlag[3]=0; refPos[4]=45; refFlag[4]=0; refPos[5]=46; refFlag[5]=0; refPos[6]=47; refFlag[6]=0; refPos[7]=48; refFlag[7]=0;  end 
14'h2256: begin refPos[0]=45; refFlag[0]=0; refPos[1]=46; refFlag[1]=0; refPos[2]=47; refFlag[2]=0; refPos[3]=48; refFlag[3]=0; refPos[4]=49; refFlag[4]=0; refPos[5]=50; refFlag[5]=0; refPos[6]=51; refFlag[6]=0; refPos[7]=52; refFlag[7]=0;  end 
14'h2257: begin refPos[0]=49; refFlag[0]=0; refPos[1]=50; refFlag[1]=0; refPos[2]=51; refFlag[2]=0; refPos[3]=52; refFlag[3]=0; refPos[4]=53; refFlag[4]=0; refPos[5]=54; refFlag[5]=0; refPos[6]=55; refFlag[6]=0; refPos[7]=56; refFlag[7]=0;  end 
14'h2260: begin refPos[0]=25; refFlag[0]=0; refPos[1]=26; refFlag[1]=0; refPos[2]=27; refFlag[2]=0; refPos[3]=28; refFlag[3]=0; refPos[4]=29; refFlag[4]=0; refPos[5]=30; refFlag[5]=0; refPos[6]=31; refFlag[6]=0; refPos[7]=32; refFlag[7]=0;  end 
14'h2261: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=35; refFlag[6]=0; refPos[7]=36; refFlag[7]=0;  end 
14'h2262: begin refPos[0]=33; refFlag[0]=0; refPos[1]=34; refFlag[1]=0; refPos[2]=35; refFlag[2]=0; refPos[3]=36; refFlag[3]=0; refPos[4]=37; refFlag[4]=0; refPos[5]=38; refFlag[5]=0; refPos[6]=39; refFlag[6]=0; refPos[7]=40; refFlag[7]=0;  end 
14'h2263: begin refPos[0]=37; refFlag[0]=0; refPos[1]=38; refFlag[1]=0; refPos[2]=39; refFlag[2]=0; refPos[3]=40; refFlag[3]=0; refPos[4]=41; refFlag[4]=0; refPos[5]=42; refFlag[5]=0; refPos[6]=43; refFlag[6]=0; refPos[7]=44; refFlag[7]=0;  end 
14'h2264: begin refPos[0]=41; refFlag[0]=0; refPos[1]=42; refFlag[1]=0; refPos[2]=43; refFlag[2]=0; refPos[3]=44; refFlag[3]=0; refPos[4]=45; refFlag[4]=0; refPos[5]=46; refFlag[5]=0; refPos[6]=47; refFlag[6]=0; refPos[7]=48; refFlag[7]=0;  end 
14'h2265: begin refPos[0]=45; refFlag[0]=0; refPos[1]=46; refFlag[1]=0; refPos[2]=47; refFlag[2]=0; refPos[3]=48; refFlag[3]=0; refPos[4]=49; refFlag[4]=0; refPos[5]=50; refFlag[5]=0; refPos[6]=51; refFlag[6]=0; refPos[7]=52; refFlag[7]=0;  end 
14'h2266: begin refPos[0]=49; refFlag[0]=0; refPos[1]=50; refFlag[1]=0; refPos[2]=51; refFlag[2]=0; refPos[3]=52; refFlag[3]=0; refPos[4]=53; refFlag[4]=0; refPos[5]=54; refFlag[5]=0; refPos[6]=55; refFlag[6]=0; refPos[7]=56; refFlag[7]=0;  end 
14'h2267: begin refPos[0]=53; refFlag[0]=0; refPos[1]=54; refFlag[1]=0; refPos[2]=55; refFlag[2]=0; refPos[3]=56; refFlag[3]=0; refPos[4]=57; refFlag[4]=0; refPos[5]=58; refFlag[5]=0; refPos[6]=59; refFlag[6]=0; refPos[7]=60; refFlag[7]=0;  end 
14'h2270: begin refPos[0]=29; refFlag[0]=0; refPos[1]=30; refFlag[1]=0; refPos[2]=31; refFlag[2]=0; refPos[3]=32; refFlag[3]=0; refPos[4]=33; refFlag[4]=0; refPos[5]=34; refFlag[5]=0; refPos[6]=35; refFlag[6]=0; refPos[7]=36; refFlag[7]=0;  end 
14'h2271: begin refPos[0]=33; refFlag[0]=0; refPos[1]=34; refFlag[1]=0; refPos[2]=35; refFlag[2]=0; refPos[3]=36; refFlag[3]=0; refPos[4]=37; refFlag[4]=0; refPos[5]=38; refFlag[5]=0; refPos[6]=39; refFlag[6]=0; refPos[7]=40; refFlag[7]=0;  end 
14'h2272: begin refPos[0]=37; refFlag[0]=0; refPos[1]=38; refFlag[1]=0; refPos[2]=39; refFlag[2]=0; refPos[3]=40; refFlag[3]=0; refPos[4]=41; refFlag[4]=0; refPos[5]=42; refFlag[5]=0; refPos[6]=43; refFlag[6]=0; refPos[7]=44; refFlag[7]=0;  end 
14'h2273: begin refPos[0]=41; refFlag[0]=0; refPos[1]=42; refFlag[1]=0; refPos[2]=43; refFlag[2]=0; refPos[3]=44; refFlag[3]=0; refPos[4]=45; refFlag[4]=0; refPos[5]=46; refFlag[5]=0; refPos[6]=47; refFlag[6]=0; refPos[7]=48; refFlag[7]=0;  end 
14'h2274: begin refPos[0]=45; refFlag[0]=0; refPos[1]=46; refFlag[1]=0; refPos[2]=47; refFlag[2]=0; refPos[3]=48; refFlag[3]=0; refPos[4]=49; refFlag[4]=0; refPos[5]=50; refFlag[5]=0; refPos[6]=51; refFlag[6]=0; refPos[7]=52; refFlag[7]=0;  end 
14'h2275: begin refPos[0]=49; refFlag[0]=0; refPos[1]=50; refFlag[1]=0; refPos[2]=51; refFlag[2]=0; refPos[3]=52; refFlag[3]=0; refPos[4]=53; refFlag[4]=0; refPos[5]=54; refFlag[5]=0; refPos[6]=55; refFlag[6]=0; refPos[7]=56; refFlag[7]=0;  end 
14'h2276: begin refPos[0]=53; refFlag[0]=0; refPos[1]=54; refFlag[1]=0; refPos[2]=55; refFlag[2]=0; refPos[3]=56; refFlag[3]=0; refPos[4]=57; refFlag[4]=0; refPos[5]=58; refFlag[5]=0; refPos[6]=59; refFlag[6]=0; refPos[7]=60; refFlag[7]=0;  end 
14'h2277: begin refPos[0]=57; refFlag[0]=0; refPos[1]=58; refFlag[1]=0; refPos[2]=59; refFlag[2]=0; refPos[3]=60; refFlag[3]=0; refPos[4]=61; refFlag[4]=0; refPos[5]=62; refFlag[5]=0; refPos[6]=63; refFlag[6]=0; refPos[7]=63; refFlag[7]=0;  end 

 default : begin refPos[0]=0; refFlag[0]=0; refPos[1]=0; refFlag[1]=0; refPos[2]=0; refFlag[2]=0; refPos[3]=0; refFlag[3]=0; refPos[4]=0; refFlag[4]=0; refPos[5]=63; refFlag[5]=0; refPos[6]=63; refFlag[6]=0; refPos[7]=63; refFlag[7]=0;  end 

endcase
 end
endmodule


